-- * IBM 360 Model 65 Emulator
-- * Copyright (C) 2024 Camiel Vanderhoeven
-- *
-- * This program is free software: you can redistribute it and/or modify
-- * it under the terms of the GNU General Public License as published by
-- * the Free Software Foundation, either version 3 of the License, or
-- * (at your option) any later version.
-- *
-- * This program is distributed in the hope that it will be useful,
-- * but WITHOUT ANY WARRANTY; without even the implied warranty of
-- * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- * GNU General Public License for more details.
-- *
-- * You should have received a copy of the GNU General Public License
-- * along with this program.  If not, see <http://www.gnu.org/licenses/>.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
USE ieee.std_logic_arith.all;


entity ROSMEM is
    Port ( clk_i : in  STD_LOGIC;
			  hclk : in STD_LOGIC;
			  rst : in STD_LOGIC;
			  hlt : in STD_LOGIC;
	        addr_i : in  STD_LOGIC_VECTOR (0 to 11);
           data_o : out  STD_LOGIC_VECTOR (0 to 99)
           );
end ROSMEM;

architecture Behavioral of ROSMEM is
  subtype ros_data_type is STD_LOGIC_VECTOR(0 to 99);
  type ros_mem_type is array(0 to 2815) of ros_data_type;
  subtype ros_address_type is integer range 0 to 2815;

  constant ros_mem_s : ros_mem_type := (
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 000
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 001
   "1000000000000000000000000100110000000000000000000111101000000011000110000000000000000000000100000000",  -- ROS word 002
   "1000001010001111000000000000111000000000000000010001001000000100000000000000000000000100010000000000",  -- ROS word 003
   "0000000000000000000010000101110000000000000000001000001101111100000010000000000000000000000100110000",  -- ROS word 080
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 081
   "1000000000000000000010000000000000000000000000001100011011111100000000000000000000000100000100000000",  -- ROS word 082
   "0000000000000000011110000011010000000000000000010110010101111100000000000010110000000100000000000000",  -- ROS word 083
   "1000000001000000000010000101111000000000000000001111100101111100000000000000000000000000000011100000",  -- ROS word 100
   "0000000000000010001010000000000000000001111000001011100110000000000010000000000000000000000100110000",  -- ROS word 101
   "1000000001000000000010000101111000000000000000001001011110000100000000000000000000000000000011100000",  -- ROS word 102
   "0000000000000000000010000101110000000000000000001100011110000100000000000000000000000000000100110000",  -- ROS word 103
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 180
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 181
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 182
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 183
   "0000000011110111100011101000001100010010100000000011000001100111001110000000000000000100000011100000",  -- ROS word 200
   "0000000011110111100011110000001100100010100000000011000001100111001110000000000000000100000011100000",  -- ROS word 201
   "0000000011110111100011111000001100110010100000000011000001100111001110000000000000000100000011100000",  -- ROS word 202
   "0000000011110111100011100000001100000010100000000011000001100111001110000000000000000100000011100000",  -- ROS word 203
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 280
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 281
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 282
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 283
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 300
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 301
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 302
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 303
   "0000000000001010000010000000000010010000000000010000011100000100000000000000000000000000000100000000",  -- ROS word 380
   "0000000000001010000000000000000101100000000100001011100010000000000000000000000000000100000100000000",  -- ROS word 381
   "0000000000000101100000000000000000000000000000001111100000000100000000000000000000000100000100000000",  -- ROS word 382
   "0000000000000000001000000000000000000000011000000110010100000000000000000000000000000100000100000000",  -- ROS word 383
   "0000001011100000000000000110011001110001100000001100000110000000000010000000000000111000000000000000",  -- ROS word 400
   "1000000000000111000000111110100000000000000011001000010011001001001111101110100000000000000100000000",  -- ROS word 401
   "1000000000000111000000111110100000000000000011001010010011001001001111001100000000000100000000000000",  -- ROS word 402
   "1000000000000111000000111110100000000000000011010010010001001001001111000100110000000000000100000000",  -- ROS word 403
   "0000000000000000000000000011011100000000000000000111100000000100000010000000000000000100000100000000",  -- ROS word 480
   "0000000110000000011100110000000111100000000000001001000100000000000001001101010100001010001000000000",  -- ROS word 481
   "0000000110000000011100110001100000000000000000010000011110000100000011001101010100001010001000000000",  -- ROS word 482
   "0000000110000000011100110000000111100000000000001001000000000000000011001101010100001010001000000000",  -- ROS word 483
   "0000001010000000000010000001001000000000000100010010001000000000000000000000000000110100010000000000",  -- ROS word 500
   "0000000000000111000010110110001000000000000000001110101001001100001111101100000000000000000100000000",  -- ROS word 501
   "0000000000000000000010000001001000000000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 502
   "0000000000000000000010000000000000000000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 503
   "1000000000000000000010000000000000000000000000001100001110000101100000000000000000000100000100000000",  -- ROS word 580
   "1000000000000111000010101110010000000000000011001011000000001100000010000000000000000100000100000000",  -- ROS word 581
   "0000000000000000000010000010100000000000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 582
   "1000000000000000000010000000000000000000000101101010100010010000000000000000000000000100000100000000",  -- ROS word 583
   "1000000000000000000010000000000000000000000110101100000000000000000010000000000000000100000100000000",  -- ROS word 600
   "1000000000000000011000000000111011000000000000101100000000000100000000000000000010000100000000000000",  -- ROS word 601
   "0000000000000000010010000000000010000000000000010000000000000110100110000000001000000100000000000000",  -- ROS word 602
   "0000000111000000011100000000000101010000000000001100000100000001101110000000000000001101110100000000",  -- ROS word 603
   "1000001011000000000000000000000000000000000000001101000000000000000010000000001010100100000000000000",  -- ROS word 680
   "0000001011001101000010000000000000000000000000001101000000000100000000000000001010000101000000000000",  -- ROS word 681
   "0000001011000000000000000000000000000000000000001101000010000001001100000000001010000001000000000000",  -- ROS word 682
   "0000000000000000010110000000000000000000000001000011101000000100000010000000000000000000000100000000",  -- ROS word 683
   "1000000001000000000000000001111000000000000000001110000000000100000000000000000000000100000011100000",  -- ROS word 700
   "1000000000000000000010000000000000000000000000001111010110000111110110000000000000000100000100000000",  -- ROS word 701
   "1000001101000100100000000000000000000000000000001110000100000100000000000000000000000000000100000000",  -- ROS word 702
   "1000000000000000001000000000000000000000000000001100100110000000000000000000000000000000000100000000",  -- ROS word 703
   "1000000000000010000010000101000000000001011000000100100110000110101100000000000000000000000001000000",  -- ROS word 780
   "0000000000000010001000000101000000000001011000010011010010000000000000000000000000000000000001000000",  -- ROS word 781
   "1000000000000010001010000101101000000001001000010011010010000000000000000000000000000000000001000000",  -- ROS word 782
   "0000000000000000000010000000000011000000000000110010100100000000000000000000000000000000000100000000",  -- ROS word 783
   "1000000010000000000000000000000000000011011000001001100010000100000000000000000000000000000100110000",  -- ROS word 800
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 801
   "0000000000000000000010000000000000000000000110100100101000000000000010000000000000000000000100000000",  -- ROS word 802
   "1000000000000100100010000000000000000000000000000101100110000100000000000000000000000100000100000000",  -- ROS word 803
   "0000000000000000000010000000000001010000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 880
   "0000000000000000000010000000000001010000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 881
   "1000000000000000000000000000000011010000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 882
   "1000000000000000000000000000000011010000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 883
   "0000000000000111000010100110000000000000000011001010100000000011000101111000100000000100000000000000",  -- ROS word 900
   "0000000000000111000010100110000000000000000011001010100100000011000101100100100000000000000100000000",  -- ROS word 901
   "1000000000100000000010000101101000000011010000010010001000000100000000000000000000000100000100000000",  -- ROS word 902
   "1000000000100000000010000101101000000011010000010010001000000100000000000000000000000100000100000000",  -- ROS word 903
   "0000001010000000000010000000000000000000000100001010010100000100000000000000000000110100010000000000",  -- ROS word 980
   "1000000000000111000010100110000000000000000011010011000000000011000101100000000000000100000100000000",  -- ROS word 981
   "1000000000000000000010000000000000000000000101101011001100010000000010000000000000000100000100000000",  -- ROS word 982
   "1000000000000000000010000000000000000000000101100000010000010000000010000000000000000100000100000000",  -- ROS word 983
   "0000000000000010000010000000000001000011011001010100000000000000000010000000000010000100000000000000",  -- ROS word a00
   "1000000000000000000010000000000000000000000110110100000000000100000000000000000000000100000100000000",  -- ROS word a01
   "1000000000010010011000000000000000000011010010010100000010000000000000000000000010000100000000000000",  -- ROS word a02
   "0000000000000010000010000000000001000011011000110100001110000000000000000000000010000100000000000000",  -- ROS word a03
   "1000000000000000000010000000000000000000000000010101000000000000000010000000000000000100000100000000",  -- ROS word a80
   "1001000000000000011110000110110000000000000000010100100000000100101111000100000000000100000100000000",  -- ROS word a81
   "0000000000000000000000000110001000000000000000010100100010000000100100000000000000000100000100000000",  -- ROS word a82
   "1000000000000111000010000110010000000000000000010101000010000000000001101100000000000100000100000000",  -- ROS word a83
   "1000001010000100100010000000000000000000000010010110000001000000000010000000000000010100010100000000",  -- ROS word b00
   "1000000000000000000000111000000000000000000100010110000010000000000000000000000000000000000100000000",  -- ROS word b01
   "1000001010000100100010000000000000000000000010110101001010000000000000000000000000000000000000001000",  -- ROS word b02
   "1000001010000000000010000000000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word b03
   "0000000000000000100000000000000000000000000011010111000010000100000010000000000000000000001000000000",  -- ROS word b80
   "0000000000000000000000000000000110010000000101110110101000000000000000000000000000000100000100000000",  -- ROS word b81
   "0000000000000000000010000000000000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word b82
   "0000000000000000000000000000000110010000000101110110101000000000000000000000000000000100000100000000",  -- ROS word b83
   "0000001011000000000000000110110000000000000000011000000010000010001000000000000000000001011000000000",  -- ROS word c00
   "0000000001000000000000000110110000000000000000011000000010000010001000000000000000000000000001000000",  -- ROS word c01
   "0000001011000000000000000110110000000000000000011000000010000010001000000000000000000000000011100000",  -- ROS word c02
   "1000000011000000000010000110110000000000000000011000000010000000000010000000000000000100000100000000",  -- ROS word c03
   "0000000000000111100010000000101000000000000000011000011111010100000001010000110000000010000111100000",  -- ROS word c80
   "0000000000000111100010000000101000000000000000011000011110000100000001010000110000000010000111100000",  -- ROS word c81
   "1000000000000111100010000100111000000000000000011000011110000100000000000000000000000000000011100000",  -- ROS word c82
   "1000000000000010000000000101101000001101001000011001000100000000000000000000000000110101011000000000",  -- ROS word c83
   "0000000000000010000000000110011000000011011000111010001110000000000000000000000000000010010010000000",  -- ROS word d00
   "1000000000000111000010000000000000001101000000011010000010000000000011001100000000000000000000000000",  -- ROS word d01
   "1000000000010000000010000010000010000011010000011101010010000000000000000000000000000100000100000000",  -- ROS word d02
   "1001011010010000000011011000000000000100001000011011101010000011111010000000000000000000110001000000",  -- ROS word d03
   "1000000000000000000010000101011000000000000000011010001000000100000010000000100000111100000100000000",  -- ROS word d80
   "1001000000000010011110000110010000000000011000010101100000000000000000000010110000000101000100000000",  -- ROS word d81
   "1000000000100111111110000000000000000101000101011000000110000000000000000010000000000100000111100000",  -- ROS word d82
   "1000000000000111111111000000000000000000000101011010000000000000000000000000100001000000000011100000",  -- ROS word d83
   "1000000000110000000010011111011000000110100100111100000000000110001000000000000000000100000100000000",  -- ROS word e00
   "0000000000000010000000000000000000001100101000011101010000000000000010000000000000000100110100110000",  -- ROS word e01
   "1000000000000010000000000000000000000000000000011100001000000100000000000000000000000000010111010000",  -- ROS word e02
   "0000000001000111000010010001000000000000000001011101010000000100000010000000000000110101011000000000",  -- ROS word e03
   "1000001011010000011110000101110000000100101000011101000000000100000011000100000000000111101101001000",  -- ROS word e80
   "1000000001010010000010000110011000000100110000011100100000000000010100000000000000000101011101000000",  -- ROS word e81
   "1000001010100000011010000000000000000100011101011101000010111100000000000000000000000000000001000000",  -- ROS word e82
   "1000001010010000000001011110000000000110010000011101000110000100000001010000100001000010000101000000",  -- ROS word e83
   "0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111",  -- ROS word f00
   "0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111",  -- ROS word f01
   "1000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000100000000",  -- ROS word f02
   "1000000000000000000010000000000000000000000000000000000000000000000000000000000000000100000100000000",  -- ROS word f03
   "0000000000001111000000000000000000001110110000011011100100000000000000000000000000000100000100000000",  -- ROS word f80
   "0000001011010000000010000000000000000101000000011111000000000100000000000000000000000100000001000000",  -- ROS word f81
   "0000001010000000011100000000000000000011011000011111000000000100000010000000100000000001000001000000",  -- ROS word f82
   "0000000000100000011100000111011000000101011100011111000010000000000000110100000000000010100000000000",  -- ROS word f83
   "0000000000000000000000000001000000000000000000000111001010000000011010000000000000000100000100000000",  -- ROS word 004
   "0000000000000010000010000001000000000011011000010001010100000100000010000000000000111100000000000000",  -- ROS word 005
   "1000000000000001000000000001000011010000000000000110101000000000011010000000000000000000000100000000",  -- ROS word 006
   "0000000000010000000010000101101000000011010000000000010110000000100100000000000000000000000100000000",  -- ROS word 007
   "1000000000000000000010000101110000000000000000001110010101111100000000000000000000000100000100110000",  -- ROS word 084
   "1000000000000000000000000101111000000000000000010111011111111100000000000000000000000000000100000000",  -- ROS word 085
   "1000000001110000000010000000000101100010100000010001010100000000000010000000000000000000000011100000",  -- ROS word 086
   "1000000001110000000010000000000101100010100000010001010100000000000010000000000000000000000011100000",  -- ROS word 087
   "0000000000000000000000000110010000000000000000010000010101111100000000000000000000000100000100000000",  -- ROS word 104
   "0000000000000010000000000001110101100000000000010001011010000000101000000000000000110000010000000000",  -- ROS word 105
   "0000000001000000000010000000000101100000000000001110011010000000000000000000000000000100000011100000",  -- ROS word 106
   "1000000000000000000010000100110101100000000000001110010010110000010110000000000000000100000100000000",  -- ROS word 107
   "0000000000000011101010000000000000000000000000001010011100000100000000000000000000000101011000000000",  -- ROS word 184
   "1000000000000010000010000000000101100000000000010001010010110000101000000000000000100100010100000000",  -- ROS word 185
   "0000000001000000000010000000000101100000000000001110011010000000110000000000000000000100000011100000",  -- ROS word 186
   "1000000000000000000010000100110101100000000000001110010010110000010110000000000000000100000100000000",  -- ROS word 187
   "1000000000000000000010000110110000000000000000000100000010000010001110000000000000000100000100000000",  -- ROS word 204
   "1000000000000000000000000010000000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 205
   "0000000001000000000010000110001000000000000000000111001000000100000000000000000000000000000100000011",  -- ROS word 206
   "0000000000000010011110000111000011010000000000001101101010000000000010000000000000000000100111100000",  -- ROS word 207
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 284
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 285
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 286
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 287
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 304
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 305
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 306
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 307
   "1000000000000010000000000011100110010011011101100111000010000000000010000000000000101101000000000000",  -- ROS word 384
   "0000000000010000000010000000000000000011010010100111001000000000011100000000000000000000000100000000",  -- ROS word 385
   "0000000100100000000000000000000000000001110000001101100100000100000000000000000000000100000100000000",  -- ROS word 386
   "1000000000000000000010000000000000000000000000000111011010000000010010000000000000000100110100000000",  -- ROS word 387
   "0000000000000111000010111110100000010000000011010000010001001001001111001000100000000100000000000000",  -- ROS word 404
   "0000000000000000000000111110100000010000000000010001000000000011010110010100100000000000000000000000",  -- ROS word 405
   "1000000000000111000010111110100000010000000011010000010001001001001111011000100000000100000100000000",  -- ROS word 406
   "0000000000000111000010111110100000010000000011010000010001001001001111010000100000000100000000000000",  -- ROS word 407
   "1000000000000000000010110000000111100000000000001001000010000000000010000000000000000100000100000000",  -- ROS word 484
   "1000000110000000000010110000000111100000000000001001000010000100000000000000000100001100000100000000",  -- ROS word 485
   "1000000110000000011100110000000111100000000000001001000000000110000000000001010100001100001000000000",  -- ROS word 486
   "0000000000000010011000000101101000000011011000000000001000000101000010000000000000000100100111100000",  -- ROS word 487
   "0000000000000000000010000000000000000000000110101010000010000100000000000000000000000000000100000000",  -- ROS word 504
   "0000000000000111000000101110010011010000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 505
   "1000000000000000000010000000000000000000000010001000010110000001100010000000000000000100000100000000",  -- ROS word 506
   "1000000000000000000000000000000011010000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 507
   "0000000000000000011110000000000010000000000000001000000110000100000000000000100000000100000000000000",  -- ROS word 584
   "1000000000010010000010000101111000000011010000001001101010010101000010000000000100000000111001000000",  -- ROS word 585
   "0000000000000111000010111110110000000000000011001011000100000011010000000000000000000000000100000000",  -- ROS word 586
   "1000000000100000000000000111000000000011010000000111101010000011001001100000000000000000000100000000",  -- ROS word 587
   "1000000000000010011110000101101101000000000000010001001100010100000001001100000000000111011111100000",  -- ROS word 604
   "1000000000000111000000000000000101000000000000001110100000000000001001001100000000000010000100000000",  -- ROS word 605
   "1000000001000111000010000101101101000000000000010000100110010100000001001100000000000111011111010000",  -- ROS word 606
   "1000000000000111000000000000000101000000000000001100000100000100001001001100000000000010000100000000",  -- ROS word 607
   "1000000000000010000000000000000000000000000000000011001000000011001100000000000000000001000110000000",  -- ROS word 684
   "0000000000000010000000000000000000000000000000000011001000000011001100000000000000000001000010010000",  -- ROS word 685
   "0000000000000010000000110000000111100000000000001001000010000000000010000000000000000101000110000000",  -- ROS word 686
   "1000000000000010000000110000000111100000000000001001000010000000000010000000000000000101000010010000",  -- ROS word 687
   "1000000000000100101000000000000000000001001000000111011110000100000010000000000000000000000100000000",  -- ROS word 704
   "1000000000001101001000000000000000000001011000010011010010000000000000000000000000000000000100000000",  -- ROS word 705
   "0000000000000000001110000000000000000000000000001011011000000100000010000000000000000000000100000000",  -- ROS word 706
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 707
   "1000000000000000000010000000000000000000000000001111000010000010001010000000000000000100000100000000",  -- ROS word 784
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 785
   "0000000101000010111110000001011000000001001000010011100100000011011011001110111010000111100000000000",  -- ROS word 786
   "1000000000000010111110000001011000000001001000010011100100000000000001001110111010000010000011110000",  -- ROS word 787
   "1000000000000000000010000000000000000000000000010000000010000100111110000000000000000100000100000000",  -- ROS word 804
   "1000000000000111100010000000000000000000000000010000011010000100000000000000000000111000000000000000",  -- ROS word 805
   "1000000000000000000010000000000000000000000000010001000110000001000100000000000000000100000100000000",  -- ROS word 806
   "1000000000000111100010000000000101110000000000000001101000000000000000000000000000111000000000000000",  -- ROS word 807
   "0000000000000000000000111110100000010000000000010001000000000011010110010100100000000000000000000000",  -- ROS word 884
   "0000000000000111100000000000000101100000000101001110010001000110001000000000000000000100110100110000",  -- ROS word 885
   "1000001010000000000000000000000010000000000100001110010001000110001000000000000000010000010100000000",  -- ROS word 886
   "0000000000000111100000000001001101100000000101001110010001000110001000000000000000000100110100110000",  -- ROS word 887
   "1000000000000110000010000101110000000000000000010011001010010101100100000000000000000100000100110000",  -- ROS word 904
   "1000000000000110000010000101110000000000000000010011001010010101100100000000000000000100110100110000",  -- ROS word 905
   "1000000000000110000010000101110000000000000000001010001110000100000000000000000000000100110100110000",  -- ROS word 906
   "1000001101000111100000000000000000000000000000010000011110000000000010000000000100000100100001000000",  -- ROS word 907
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 984
   "1000000011000000000010000001111000000000000000010010001010000000000000000000000000000100000100000000",  -- ROS word 985
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 986
   "0000000011000000000010000001111000000000000101100000000110010000000010000000000000000000000100000000",  -- ROS word 987
   "1000000000000000001000000000000000000000000000110100000000000100000010000000000000000000000100000000",  -- ROS word a04
   "0000000000000000000010000000000011110000000000010100000010000100000010000000000000000000000100000000",  -- ROS word a05
   "0000000000000000000010000000000000000000000010010100000010000001100010000000000000000000000100000000",  -- ROS word a06
   "1000000000000000000010000000000000000000000110110100000100000000000000000000000000000100000100000000",  -- ROS word a07
   "0000000000000111000000000110011000000000000000010100100010000100000011001100000000000110000100000000",  -- ROS word a84
   "1000000000000000011100000000000000000000011000010100100100000000000000000010000000000100000000000000",  -- ROS word a85
   "0000000000000000000010000000000000000000000001010101000010000100000010000000000000000000000100000000",  -- ROS word a86
   "1011010000100000000000000000000000001000011001010101000100000000000000000000000000000000000100000000",  -- ROS word a87
   "0000000000000111100010000000000000000000000000010110000010000100000000000000000000000000110100110000",  -- ROS word b04
   "0000000000000000000000111000000000000000000010010110001000000010100010000000000000000100000100000000",  -- ROS word b05
   "0000000000000000000000111000000000000000000101010110000001000000000000000000000000000100000100000000",  -- ROS word b06
   "1000001010000000000010000000000000000000000010110101001010000000000000000000000000000000000000001000",  -- ROS word b07
   "1000000000000111000000000110110000000000000000010110100110000100000011001100000000000100000000000000",  -- ROS word b84
   "0000000000000111000000000000000010100000000000010110101010000100000011001111110000000110000100000000",  -- ROS word b85
   "0000000000000000000000000000000110010000000101101111000110000100000000000000000000000100000100000000",  -- ROS word b86
   "0000000000000000000010000110110000000000000011110111000010000100000000000000000000000000000100000000",  -- ROS word b87
   "1000001001010111100000000100101000000101010101011000001010000000000000010000000000000100110000110000",  -- ROS word c04
   "0000001001010111100010000100101011010101010101011000001010000000000000010000000000000100110000110000",  -- ROS word c05
   "0000000000000000011100000000000000000000000000011000001010000000000010000000100000000000000000000000",  -- ROS word c06
   "0000000000000000000010000101011000000000000101011000010110000010001001110100000000111010000100000000",  -- ROS word c07
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word c84
   "0000000000010111000000000110011000000011010000011001000100000001100101101110100000000010000000000000",  -- ROS word c85
   "1000000000001111000000000001000001010000000000011001100000000000001100000000000000010100000000000000",  -- ROS word c86
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word c87
   "0000000000000111100000000100101000000000000000011010000010000100000100000000000000000100110100110000",  -- ROS word d04
   "1000000000010000000010000000000000000011010000011010001100000000000010000000000000000100000100000000",  -- ROS word d05
   "0000000000001111000010000001001000000000000000011010000100000000000000000000000000000101011000000000",  -- ROS word d06
   "0000001010000010000000000110101000001101010000011010101010000000000000000000000000111100010100000000",  -- ROS word d07
   "0000000000000111000000000101011000000000000000011011000010000100000011001100000000000011101001001000",  -- ROS word d84
   "0000000000000111000000000101011000000000000000011011000010000100000010000000000000000001101001001000",  -- ROS word d85
   "1000001010000111000010011110011000001110101100111011100010000000000011010000100000000010000001000000",  -- ROS word d86
   "0011110000000010000000000000000000000000000000011011000100000000000000000000000000000001011000000000",  -- ROS word d87
   "0000001010000000000010000010111000000000000100011101011100000100000000000000000000010000010100101000",  -- ROS word e04
   "1000001010000000000010000010111000000000000100111100000010000100000010000000000000010100010100101000",  -- ROS word e05
   "1000001010000000000000010010111000000000000100011101011000000100000010000000000000000001000111100000",  -- ROS word e06
   "1000000000000010000000011000000000001100101000011100001010000000000000000000000000000000000100110000",  -- ROS word e07
   "0000000000000000000010000000000000000000000000011101000010000100000010000000000000000000000100000000",  -- ROS word e84
   "1000000001000010000010000000000000001100101010011101010000000000000000000000000000000100110100110000",  -- ROS word e85
   "0000000000000000011010000000000000000000000000011101000010000100000010000011110000000000000100000000",  -- ROS word e86
   "0000000000010111100010000000000000000100000100111101001010000100000001000100000000000010000111100000",  -- ROS word e87
   "0000000000001111010110100101101000001110000000011110000100100010001001010000100001000110000000000000",  -- ROS word f04
   "1000000000000010010100001110011000001100010000011101010100000100000010000000100001000100010000000000",  -- ROS word f05
   "0000001010000000000010000010111000000000000011011110000111011000011010000000000000000100010001001000",  -- ROS word f06
   "1000001011000000000000000000000000000000000101011110001010000100000010000000000000000101101000110000",  -- ROS word f07
   "0000001101011111000010000000000000000100111000011111000010000100010100000000000000000000000100000000",  -- ROS word f84
   "1000000000010010000000000101011000000110001000011111001010000100000010000000000000000000001111100000",  -- ROS word f85
   "0000000000010111100000000101110000000100010000011101000001011100000001101100000000000110000101000000",  -- ROS word f86
   "1000000000000111000010000110110000001101011000011111000100000000000110000000000000000100000100000000",  -- ROS word f87
   "1000000000000001000000000001000011010000000000000110101000000000011010000000000000000000000100000000",  -- ROS word 008
   "0000000000000000010100000101001000000000000110110010010100000000100110000000000000000100000100000000",  -- ROS word 009
   "0000000000000001000000000001000011010000000010000110101000000000011010000000000000000100000100000000",  -- ROS word 00a
   "1000000000001011011100011000111000000000000000000000010100000100000010000000000000111100000000000000",  -- ROS word 00b
   "0000000110000000000011001000000000000000000000000110100000000011110100000000000000000100000011100000",  -- ROS word 088
   "0000000110000000000011001000000000000000000000000101100000000011110100000000000000000100000011100000",  -- ROS word 089
   "1000000110000000000011001000011000000000000000000110100000000011110100000000000000001100000111100000",  -- ROS word 08a
   "0000000110000000000001001000010000000000000000000101100000000011110100000000000000001100000111100000",  -- ROS word 08b
   "1000001011000000000000000000000000000000000000001111100001111100000000000000001010100100000000000000",  -- ROS word 108
   "1000000001000000000000000000000000000000000000001101000001111100000000000000000000000100000011100000",  -- ROS word 109
   "1000000001000000000000000000000000000000000000001101000001111100000000000000000000000100000011100000",  -- ROS word 10a
   "1000000001000000000000000000000000000000000000001101000001111100000000000000000000000100000011100000",  -- ROS word 10b
   "1000001011000000000000000110000000000000000000001001011100000100000000000000000000000100000001000000",  -- ROS word 188
   "0000001011000000000010000110111000000000000000001111011100000100000000000000000000000100000001000000",  -- ROS word 189
   "0000000000000000000010000010100000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 18a
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 18b
   "1000000000000010000000000000000000000000000000000100010100010100000000000000000000000000000100110011",  -- ROS word 208
   "1000000000010000000001111011000000000000110000000100000100101000000000000000000000000100010010100000",  -- ROS word 209
   "0000000000000011100000000000000000000000000000000100010100010100000000000000000000000000000000110010",  -- ROS word 20a
   "1000000000000000000010000000110000000000000000000100010100000000000010000000000000000100000100000000",  -- ROS word 20b
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 288
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 289
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 28a
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 28b
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 308
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 309
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 30a
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 30b
   "1000000000000000000000000001000011000000000110101101011000000100000000000000000000000000000100000000",  -- ROS word 388
   "1000000000110111100010000000001000000001110101000010000000000011001110000000000000000101011111100000",  -- ROS word 389
   "0000000000000000000010000000000000000000000000000110000000000011001110000000000000000000000100000000",  -- ROS word 38a
   "0000000000000000000010000000000000000000000000001000011000000011001100000000000000000000000100000000",  -- ROS word 38b
   "1000000000000111111100000000000000000000000000010001100110011001000011111100000000000010110100110000",  -- ROS word 408
   "0000000000001101000000000000000000000001111000101000001000000000000010000000000000000100000100000000",  -- ROS word 409
   "1000000000000000000010000000000000000000000000010011000110000000101010000000000000000100000100000000",  -- ROS word 40a
   "1000000000000000000010000000000000000000000000010000001110000100000010000000000000000100000100000000",  -- ROS word 40b
   "1000000110000111011100110110010111100000000000001001000010000100000001001101010100001110001000000000",  -- ROS word 488
   "1000000000000010000010000000000110010011011101001111010100000100000000000000000000000001000000000000",  -- ROS word 489
   "0000000000000010000000000000000000000001111000001011100110000000000010000000000000000000000001000000",  -- ROS word 48a
   "1000000000000010000010000000000000000001101000001011100110000000000010000000000000000000000001000000",  -- ROS word 48b
   "0000001010000000000010000001001000000000000100010010001000000000000000000000000000110100010000000000",  -- ROS word 508
   "1000000000000111000010110110001000000000000000001111101001001100001111101100000000000100000100000000",  -- ROS word 509
   "0000000000000000000010000001001000000000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 50a
   "0000000000000000000010000000000000000000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 50b
   "0000000000000111100010000111100000000000000000001011000010000100000000000000000000011000000100110000",  -- ROS word 588
   "0000001011000000000000000110011000000000000000001101010000000100001110000000000000011100000100000011",  -- ROS word 589
   "0000000000000000000010000000000000000000000101101011000000101100000000000000000000000000000100000000",  -- ROS word 58a
   "0000001011000000000000000110011000000000000000001101010000000100001110000000000000011100000100000011",  -- ROS word 58b
   "0000000110000000011110010000000101000000000000010000100100000100100011001100000000001110101000000000",  -- ROS word 608
   "1000000110000000011110010000000101000000000000010000100100000000100011001100000000001010101000000000",  -- ROS word 609
   "1000000000000010000000000000000000000001111000001110100010010100000000000000000000000001011111010000",  -- ROS word 60a
   "0000000000000010000000000000000000000001111000001110100010010100000000000000000000000001011000000000",  -- ROS word 60b
   "1000000000000111100010000000000000000000000000001111000100000000000010000000000000000100110100110000",  -- ROS word 688
   "0000000011000000000000000000010000000000000000001101000110000100000110000000000000000100000100000000",  -- ROS word 689
   "0000001010000000000010000000000000000000000100001101010100000100000000000000000000010000010100000000",  -- ROS word 68a
   "0000000000100000000010000000000000000011010000010001011000000000000010000000000000000000000100000000",  -- ROS word 68b
   "0000000000000000000010000000000000000000000000001110000010000000101100000000000000000000000100000000",  -- ROS word 708
   "0000000000000000011100000000000000000000000000000111100000000011110001001100000000000110000100000000",  -- ROS word 709
   "0000000000000111111100000000110000000000000000001110000100100000000010011101100000000100000101000000",  -- ROS word 70a
   "1000000000000000011100000101101000000000000000000001100000000011110111001110000000000110000000000000",  -- ROS word 70b
   "1000000101000000000000000110100101000000000000000100100110000000111000000000000000000000101101010000",  -- ROS word 788
   "0000001010000000000010000110010101100000000100001111000100000100000000000000000000010000010100000000",  -- ROS word 789
   "1000000000000000000010000110110000000000000000001111001110000100101110000000000100000100010110100000",  -- ROS word 78a
   "1000000000000111100010000000000000000000000001101010000100000000000000000000000000000000000000100000",  -- ROS word 78b
   "1000000110000000000011001000000000000000000000000110100000000011000000000000000000000000000011100000",  -- ROS word 808
   "1000000110000000000011001000000000000000000000000101100000000011000000000000000000000000000011100000",  -- ROS word 809
   "0000000110000000000011001000011000000000000000000110100000000011000000000000000000001000000111100000",  -- ROS word 80a
   "1000000110000000000001001000010000000000000000000101100000000011000000000000000000001000000111100000",  -- ROS word 80b
   "0000000000000000000010011000000000000000000010010000011100000100000000000000000000000101000000000000",  -- ROS word 888
   "1000000000000000000010011000000000000000000011010000011100000100000000000000000000000001000000000000",  -- ROS word 889
   "0000000000000000000010000011010110010000000101110001000100000001001010000000000100000000010110100000",  -- ROS word 88a
   "0000000000000000000000011000000000000010011000010000011100000100000000000000000000000001000000000000",  -- ROS word 88b
   "1000000100010000011110000000000000000011010000010010000010000100000011001111000000011010011001110000",  -- ROS word 908
   "0000000100010000011110000000000000000011010000010010000010000100000011001101000000011010011101110000",  -- ROS word 909
   "1000000000000110000000110110001000000000000000001010101001001100001111110100000000000100000000100000",  -- ROS word 90a
   "1000000000000110000000101110010000000000000011001011000000001100000010000000000000000100000000100000",  -- ROS word 90b
   "0000001001000000000010000000000000000000000000001001100100000000000010000000000000000000000100000000",  -- ROS word 988
   "0000000001000000000000000000000000000000000000001001100100000000000010011110110000000000000011100000",  -- ROS word 989
   "0000001001000000000010000000000000000000000000001001100100000000000010000000000000000000000100000000",  -- ROS word 98a
   "0000001001000100100010000000000000000000000000001001100100000000000010011110110000000000000100000000",  -- ROS word 98b
   "1000000000000000000010000000000000000000000000010100000100000000000010000000000000000100000100000000",  -- ROS word a08
   "1000001001000000000000000000000010110000000001010100000100000100000000000000000000000000000100000000",  -- ROS word a09
   "1000000000000000000010000000000000000000000001010100000100000100000010000000000000000100000100000000",  -- ROS word a0a
   "1000000000000010000010000000000001000011011000110100000110000000000000000000000010000000000000000000",  -- ROS word a0b
   "1000000000000000000010000000000000000000000000010101000100000000000010000000000000000000000011100000",  -- ROS word a88
   "0000000000000010000000000000000000000000000000010100100100000100010100000000000000000001000000000000",  -- ROS word a89
   "1000000000000000000010000110011000000000000001010101000110000000000000000000000000000100000100000000",  -- ROS word a8a
   "0000000000000000000000000110011000000011111001010101000110000000000000000000000000000100000100000000",  -- ROS word a8b
   "0000000000000111100000111000000000000000000101010111100001000000000000000000000000000100110100110000",  -- ROS word b08
   "0000000000000000000010000000000000000000000100010111101000000000000000000000000000000000000100000000",  -- ROS word b09
   "1000001010000000000010000000000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word b0a
   "1000001010000000000010000000000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word b0b
   "0000000000000000000010000001111000000000000000010001010110000000111100000000000000000000000100000000",  -- ROS word b88
   "1000000000000011100000000000000000000011011000010111000110000000000000000000000000111100000000000000",  -- ROS word b89
   "1000000000000111100010000000000000000000000000010001001000000100011010000000000000110000010000000000",  -- ROS word b8a
   "1000000000000000000010000001001010100000000000010101001110000100000010000000000000000100000100000000",  -- ROS word b8b
   "0000000000100000010110010000000000000010001000011000011010000100000000000010000000000100000000000000",  -- ROS word c08
   "0000000000000010011110000000000000001101010000011000010100000110001010000010000000111101011000000000",  -- ROS word c09
   "1000000000000000010110000101110000000000000000011000001000001110100010000000000000011100000100000000",  -- ROS word c0a
   "0000000001110000000000000110011000000101000000011000011100000000000010000000000000000100110100110000",  -- ROS word c0b
   "1000000000010111100010000000000000000011010101011001000100000100000010000000000000000100110100110000",  -- ROS word c88
   "0000000000000111100000000000000000001101000101011001000100000100000010000000000000000100110100110000",  -- ROS word c89
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word c8a
   "1000001001000010000000000000000000000000000010011000011100000000000000000000000000000100000000001000",  -- ROS word c8b
   "0000000000000010000000000000000000001101010000011010000110000100000000000000000000111100010100000000",  -- ROS word d08
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d09
   "0000000000010000000010011110110000000011010000011010001010000110001010000000000000000000000100000000",  -- ROS word d0a
   "1000000000010000000010000110110000000011010000011010000000000000000010000000000000000100000100000000",  -- ROS word d0b
   "1000000001010111000010000110100000000100001000011011000100000000000011001100000000000100000101000000",  -- ROS word d88
   "0000001011000111000010000000000000000000000000011011000100000100000001001100000000000101011000111000",  -- ROS word d89
   "0011110000010010000010010110000000000100101000011010000110000000000010000000000000000100000001000000",  -- ROS word d8a
   "0000000000000000000010000000000000000000000000010101100110000000000010000000000000000000000100000000",  -- ROS word d8b
   "0000000001000000000000000000000000000000000111011100001000000100000010000000000000110001011000000000",  -- ROS word e08
   "0000001011001111010101010000000000000000000000011101001111010100000010000010100001110000000000000000",  -- ROS word e09
   "1000000000100000000010000000011000000110100100111100000110000010001000000000000000010000000000000000",  -- ROS word e0a
   "0000000001000111100000000000000000000000000111011100000110000110001010000000000000000100110100110000",  -- ROS word e0b
   "1001010000001010000000000000000010000000000001011101001000000000000010000000000000000000000100000000",  -- ROS word e88
   "0001010000101010010100100000000000000100011001011101000110000000000011010000100001000100000100000000",  -- ROS word e89
   "1001010000001010010100100000000000000000000001011101000110000000000001010000100001000000000100000000",  -- ROS word e8a
   "1000000000000000010110101000000000000000000000011101000110000100000011010000100001000100000100000000",  -- ROS word e8b
   "0010100000000111000000000110110000000000000011011110000010000100000000000000100001000100000100000000",  -- ROS word f08
   "0000000000000000011100000110011000000000000101011110011100000110001011000100000000000010000000000000",  -- ROS word f09
   "1010100000000111000010000110110010000000000011011110000010000100000000000000100001000100000100000000",  -- ROS word f0a
   "0000000000000000000010000000000000000000000101011110010010000110001011000100000000000110000000000000",  -- ROS word f0b
   "1000001001000011100010000110110000001100111000011111000100000100000010000000000000000101000101011000",  -- ROS word f88
   "0000000000000111100010000101110000000000000101011100010010000110001000000000000000000100000001000000",  -- ROS word f89
   "1000000000000010011100000110010000001100110101011111000110000100000010000000000000000001011111100000",  -- ROS word f8a
   "1000000000010010000000000001110000000100010000011111000110000000000000000000000000000000000100000000",  -- ROS word f8b
   "0000000000000001000010000001000001010000000000000110101000000000011010000000000000000000000100000000",  -- ROS word 00c
   "1000000000000111111010000000000000000000000000110001101010001001001111001111110000000010110000100000",  -- ROS word 00d
   "1000000000000000000010000001000011010000000000010010100010000100011010000000000000000100000100000000",  -- ROS word 00e
   "1000000000000000000010000100100000000000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 00f
   "0000000011010000000001001000000000000001100000001100100001111111110100000000000000000000000011100000",  -- ROS word 08c
   "0000000011110000000011001000000000000001100000001101100001111111110100000000000000000100000011100000",  -- ROS word 08d
   "0000000011010000000001001000011000000001100000001100100001111111110100000000000000000000000011100000",  -- ROS word 08e
   "1000000011110000000001001000010000000001100000001101100001111111110100000000000000000100000011100000",  -- ROS word 08f
   "1000001011000000000001000110111000000000000000001101000111111100000000000000001010100100000000000000",  -- ROS word 10c
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 10d
   "0000000000000000000000000011010000000000000000001101000101111100000010000000000100000100010110100000",  -- ROS word 10e
   "0000000000000000000010000110011000000000000000010010000111111100000000000000000000000000000100000000",  -- ROS word 10f
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 18c
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 18d
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 18e
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 18f
   "0000000000000010000000000000000000000000000000000100010110010100000000000000000000000100000100110011",  -- ROS word 20c
   "1000000000010000000010000011000000000000111000000100000110101000000000000000000000000000010010100000",  -- ROS word 20d
   "1000000000000011100000000000000000000000000000000100010110010100000000000000000000000100000000110010",  -- ROS word 20e
   "1000000000000000011110000110111000000000000000001100001000000011001100000000100000000000000000000000",  -- ROS word 20f
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 28c
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 28d
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 28e
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 28f
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 30c
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 30d
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 30e
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 30f
   "1000000000001010000010000011000000000000000000100100011100101000000000000000000000000000010010100000",  -- ROS word 38c
   "0000000000000000000001110011000000000000000000000100011110101000000000000000000000000000010010100000",  -- ROS word 38d
   "0000000000000010000011101000000000000011011000000111011000010100000000000000000000010000010100000000",  -- ROS word 38e
   "1000000000000010000011101000000000000011011000000111011000010100000000000000000000000000010000000000",  -- ROS word 38f
   "1000000001000000011100000110111000000000000000001100010000000000000000000000100000000000000111100000",  -- ROS word 40c
   "0000000000000111000000000000000000000000000000001011010000000000000011001100000000000000000000000000",  -- ROS word 40d
   "0000000000000000000010000111100000000000000000001011000010100000000000000000000000000000000100000000",  -- ROS word 40e
   "0000000000000000000010000111100000000000000000001011000010100000000000000000000000000000000100000000",  -- ROS word 40f
   "0000000000010010000001000000000000000001100000001110100100000100000010000000000000000000000001000000",  -- ROS word 48c
   "1000000000010010000000000001001000000011010000001001000110000100001000000000000000000101011000000000",  -- ROS word 48d
   "0000000110100000000011000000000000000010100000001110100100000100000010000000000000000001000111010000",  -- ROS word 48e
   "1000000110100000000011000000000000000010100000001110100100000100000010000000000000000000000011010000",  -- ROS word 48f
   "1000000000000111100010000000000000000000000101001010000110000100000000000000000000000000000000100000",  -- ROS word 50c
   "0000000000000111000000101110010011010000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 50d
   "0000000000000010000000000000000000000000000000100010101010000100000010000000000000000001011000000000",  -- ROS word 50e
   "1000000000000000000000000000000011010000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 50f
   "1000000000000111100010000000000000000000000000010000011000000000001110000000000000011100000100110000",  -- ROS word 58c
   "1000001011000000000000000110011000000000000000001101010000000000001110000000000000011000000100000011",  -- ROS word 58d
   "0000000000000000000010000001001000000000000101101011000000101100000000000000000000000000000100000000",  -- ROS word 58e
   "1000001011000000000000000110011000000000000000001101010000000000001110000000000000011000000100000011",  -- ROS word 58f
   "1000000110000000000010000000000101000000000000001100000000000100000010000000000000001100101100010000",  -- ROS word 60c
   "0000001101000010000010000000000000000011011000001001000110000001100100000000000000001000000111010000",  -- ROS word 60d
   "0000000110000000000010000000000101000000000000001100000000000100000010000000000000001100101001100000",  -- ROS word 60e
   "0000000000010010000000000000000000000011010000010010000110000000000010000000000000000000000001000000",  -- ROS word 60f
   "0000001011000000000000000000000000000000000000001110011110000100000010000000001010000001000000000000",  -- ROS word 68c
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 68d
   "0000000000001100011100000001111000000011011000010010011110000000000010000000101010000000000000110000",  -- ROS word 68e
   "0000000000000010000000000000000000000011011000000000011110000100000000000000000000000000000011010000",  -- ROS word 68f
   "0000000000000000000010000000000000000000000110101110011000000100000000000000000000000000000100000000",  -- ROS word 70c
   "0000000001000000000010000001111010000000000000001110000000000100000000000000000000000100000011100000",  -- ROS word 70d
   "0000000000000000000010000011101000000000000000001110100110000100010100000000000000000000000100000000",  -- ROS word 70e
   "1000000011110000000010000001001000001000010000010111010100000000000000000000000000000100000100000000",  -- ROS word 70f
   "0000000000000000000000000000000000000001011000010011100110000000000000000000000000000100000100000000",  -- ROS word 78c
   "0000000000100111111100000000000000000011010000010001100100000000010010000000100000000100000100100000",  -- ROS word 78d
   "0000000110000000000010000101101101110000000011000110101000000100000010000000000000010100110000000000",  -- ROS word 78e
   "0000000000000111000010000001011000000001001000010011100100000000000001001100100000000000000100000000",  -- ROS word 78f
   "1000000011010000000001001000000000000001100000001100100001111111000000000000000000000100000011100000",  -- ROS word 80c
   "1000000011110000000011001000000000000001100000001101100001111111000000000000000000000000000011100000",  -- ROS word 80d
   "1000000011010000000001001000011000000001100000001100100001111111000000000000000000000100000011100000",  -- ROS word 80e
   "0000000011110000000001001000010000000001100000001101100001111111000000000000000000000000000011100000",  -- ROS word 80f
   "0000000000000000000010000000000000000000000000010001001000000010101010000000000000000000000100000000",  -- ROS word 88c
   "0000000000000000000000000101100000000000000000001000100000000100000010000000000000000100000100000000",  -- ROS word 88d
   "0000000000000000000010000000000000000000000000010000000010000000110010000000000000000000000100000000",  -- ROS word 88e
   "1000000000000011100000000000000000000011011000010001011010000100000000000000000000111100000000000000",  -- ROS word 88f
   "0000001011000100100000000000000000000011011000101010011110000000000010000000000000000100000100000000",  -- ROS word 90c
   "1000000000000000000010011000000000000011011000001000100100000100000010000000001010000001001000000001",  -- ROS word 90d
   "0000000000000000000010000101101000000000000000010010101000000100000000000000000000000000000100000000",  -- ROS word 90e
   "1000000110000010100010000000000000000000000000001001011110000000000011100000000000000010100001110000",  -- ROS word 90f
   "0000000000000000000010000000000000000000000000001000000100000101000100000000000000000000000100000000",  -- ROS word 98c
   "1000000000000010000000000000000000000000000000000000011110000100000010000000000000111100000000000000",  -- ROS word 98d
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 98e
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 98f
   "0000000000010010000010000000000000010011010000110100000110000000000010000000000010000100000000000000",  -- ROS word a0c
   "0000000000000000000010000000000011110000000000010100000110000100000000000000000000000000000100000000",  -- ROS word a0d
   "0000000000000000000010000000000000000000000110110100000110000100000010000000000000000000000100000000",  -- ROS word a0e
   "1000000000000000000010000000000000000000000010010100001000000000000000000000000000000100000100000000",  -- ROS word a0f
   "0000001011000000000000000110010000000000001000110101000110000100000000000000000000100000000000000000",  -- ROS word a8c
   "0000000000000010011110000000000000000000000000010101001000000000000010111100110000000011011100000000",  -- ROS word a8d
   "0000001011000000000000000011101000000000000001010101000110000100010100000000000000011001000000000000",  -- ROS word a8e
   "1000000000000000000010000011110000000000000000010101100010000000000010000000000000000100000100000000",  -- ROS word a8f
   "1000000000000000000010000000000000000000000100010110001000000100000000000000000000000100000100000000",  -- ROS word b0c
   "1000000000000000000000111000000000000000000101010110010010000000000000000000000000000000000100000000",  -- ROS word b0d
   "0000000000000000000010000000000000000000000101010110001010000100000010000000000000000000000100000000",  -- ROS word b0e
   "0000000000000000000010000000000000000000000101010110001010000100000010000000000000000000000100000000",  -- ROS word b0f
   "0000000000010000000010000000000000000011010000010111000110000000000010000000000000000000000100000000",  -- ROS word b8c
   "0000000000001001000010000000000000000000000000010111000110000100000000000000000000000000000100000000",  -- ROS word b8d
   "0000000000000000000000000000000000000000001000010111000110000100000010000000000000000100000100000000",  -- ROS word b8e
   "0010010000000000011100000000000000000000000000010000011100000100000000000010110000000000000000000000",  -- ROS word b8f
   "1000000000011111000000000100000000000101010000011000000110000000000010000000000000000000000100110000",  -- ROS word c0c
   "0000000000100111100010000000000000010101101101011000000110000100000001010010100000000010000111100000",  -- ROS word c0d
   "0000001001010000000001000110011000000101100010011000001100001100000000000000000000000000000001000000",  -- ROS word c0e
   "1000000000000010000010000111101000000011011000011000001110000110001001001000100000000101000100000000",  -- ROS word c0f
   "1000000000000010000010000000000000001101101000011001000010100000000000000000000000000001011000000000",  -- ROS word c8c
   "1000000000000010000010000100001000001101101000011001000010100000000000000000000000000001011000000000",  -- ROS word c8d
   "1000000000100000010110000111011000000101000101011001000010000000000010000010000000000000000000000000",  -- ROS word c8e
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word c8f
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d0c
   "1000000000000110000010010110100000000000000000011010001110000100000011001100000000000100000101000000",  -- ROS word d0d
   "1000001010100000000000000000000000000110000000011010010000000000000010000000000000000000000100110000",  -- ROS word d0e
   "0000000001000000000000000000000000000000000000011011010010000000000010000000000000110001011000000000",  -- ROS word d0f
   "0000000000000010000010000000000111000000000000010101100010000100000010000000000000000000000100000000",  -- ROS word d8c
   "1000000000000000000000000110010000000000000000010100011101111100000010000000000000000000000100000000",  -- ROS word d8d
   "1010001011010000000010000000000000001000000000010111001110000100000000000000000000000100000100000011",  -- ROS word d8e
   "0000000000010010000010000110011000000100111000011111000000000000000010000000000000000100010000000000",  -- ROS word d8f
   "1000000001000000000010000001000000000000000001011101010000000100000010000000000000000101011111010000",  -- ROS word e0c
   "1000000000000000000010110000000000000000000000011101001100000110001010000000000000000100000100000000",  -- ROS word e0d
   "1000000000000010000000000000000000001100101010011101001000000110000100000000000000000000110100110000",  -- ROS word e0e
   "1000001011001111010111110000000001010000000000011101001111010100000010000010100001110000000000000000",  -- ROS word e0f
   "0000000001001011110110001110110000000000000000011110001110000000000001010000100001000010000100001000",  -- ROS word e8c
   "0000000000011011100000000000000000000100111000011110010100000010001000000000000000000100000100000000",  -- ROS word e8d
   "0000000000111111000010000000000000000100100000011100001000000010001000000000000000000100000001000000",  -- ROS word e8e
   "0000000000001111011010000110011000000000000000011101001010000000000000000000000000000100000011100000",  -- ROS word e8f
   "0000001011000000000000000000000000000000000000011110001000000000011110000000000000000001101000110000",  -- ROS word f0c
   "1000000000000000000010000000000000000000000100111110001000000100011110000000000000000100000100000000",  -- ROS word f0d
   "1000001011000000000010111000000000000000000000011110001000000000011110000000000000000001101000110000",  -- ROS word f0e
   "0000000000000000000000111000000000000000000100111110001000000100011110000000000000000100000100000000",  -- ROS word f0f
   "1000001010000111000010000110100000000000000100111111000110000000000011001100000000000100000101000000",  -- ROS word f8c
   "1000000000000111000000000101110000001101001000011111000110000100000001001100000000000100000000110000",  -- ROS word f8d
   "0000000001100000000000000110011000000101010000011111000100000100000000000000000000000000000011100000",  -- ROS word f8e
   "1001010000101010011010111000000000000100100000011111001000000100000010000011100001000100000100000000",  -- ROS word f8f
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 010
   "0000000000000000010100000101001000000000000110101101000000000100000010000000000000000100000100000000",  -- ROS word 011
   "0000000000010010000000000111000011010011010000001101101010000000000010000000001010000001001001000000",  -- ROS word 012
   "0000000000010010000010000111000000000011010000001111001010000000000000000000001010000101001001000000",  -- ROS word 013
   "1000000000000000000010000000000000000000000000001000001011111100000000000000000000000100000100000000",  -- ROS word 090
   "1000000001000000000010000101111000000000000000001001011100000000000010000000000000000100000100000011",  -- ROS word 091
   "0000000001000000000010000101111000000000000000010001011100000000000000000000000000000000000100000011",  -- ROS word 092
   "1000000000000000000000000101110111110000000000010001011010000100000010000000000000000000000100110000",  -- ROS word 093
   "1000000000000000000000000011010000000000000011101011100111111100000010000000000100000000010110100000",  -- ROS word 110
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 111
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 112
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 113
   "0000000000000000000010000000011000000000000000010010011110000100000010000000000000000100000011100000",  -- ROS word 190
   "0000000000000000000010000000011000000000000000010001011110000100000010000000000000000100000011100000",  -- ROS word 191
   "0000000000000000001000000000011000000001111000001001001010000000000010000000000000000000000011100000",  -- ROS word 192
   "1000000000000010001010000000011000110001111000001001001010000000000010000000000000000000000011010000",  -- ROS word 193
   "1000000001100000000001110000000100100010100000000111000101100100000010000000000000000100000011100110",  -- ROS word 210
   "1000000001100000000001111000000100110010100000000111000101100100000010000000000000000100000011100101",  -- ROS word 211
   "0000000001100000000000000000000100000010100000000111000101100100000010000000000000000100000111100100",  -- ROS word 212
   "0000000001100000000001101000000100010010100000000111000101100100000010000000000000000100000111100111",  -- ROS word 213
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 290
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 291
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 292
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 293
   "1000000000001111011000000000000011100000000000110000100010000100000010000000000010000100000000000000",  -- ROS word 310
   "0000000000000111000000000000000000000000000000001001010110000110001111101110100000000100000100000000",  -- ROS word 311
   "0000000000000111000000000000000000000000000000001011010110000110001111001100000000000000000000000000",  -- ROS word 312
   "1000000000000111000000000000000000000000000000001000010110000110001111000100110000000000000100000000",  -- ROS word 313
   "0000000000000000000010000010001000000000000000010110100110000010100010000000000000000000000100000000",  -- ROS word 390
   "0000000000000010000000000000000000000000000000010110100110000010100010000000000000000000000000001000",  -- ROS word 391
   "0000001010000000011100000000000000000000000000000110011010000010100101001100000000110100010100000000",  -- ROS word 392
   "1000000000000010000000000000000000000011011000000111001110010100000000000000000000000100010000000000",  -- ROS word 393
   "0000000000010111100000001000000000000001110101000110001100000001000010000000000000000100110100110000",  -- ROS word 410
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 411
   "1000000001010000011010000111000000000011010000010000101010000011001000000011000100000000111011100000",  -- ROS word 412
   "0000000001010000011010000111000000000011010000010000101010000011001000000001000100000000111111100000",  -- ROS word 413
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 490
   "0000000000000010000000000000000000110001111000001001001000000000000000000000000000000000000011010000",  -- ROS word 491
   "1000000000000000000000011000000010000000000000001000001000000110101000110100000000000110000001000011",  -- ROS word 492
   "0000000000000000000010011101101000000000000000001000001000000110101000110100000000000110000001000011",  -- ROS word 493
   "0000000001000000000000000000000000000000000000001010001110000000000010000000000000000100101100000000",  -- ROS word 510
   "1000000000000000000000000000000001110000000000000110011100000000010100000000000000000000000100110000",  -- ROS word 511
   "0000000000000010001010000000100000000001101000001001001000000000000000000000000000000000101100000000",  -- ROS word 512
   "0000000000000111000000110110000000000000000000010001001011001100001111101000001000000100000100000000",  -- ROS word 513
   "0000000000000000000010000000000000000000000000001110011110000000000000000000000000000000000100000000",  -- ROS word 590
   "0000000000000010000010000000000001000011011000101011001000000100000000000000000010000100000000000000",  -- ROS word 591
   "0000000000010010000010000000000000010011010000101010000010000000000000000000000010000100000000000000",  -- ROS word 592
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 593
   "0000000000000111000010000110010000000000000000001011010000000100000000000000000000000000000100000000",  -- ROS word 610
   "1000000000000111100000000000000010000000000000010010000000101110101000000000000000000100000000100000",  -- ROS word 611
   "0000000000000111000000000000000000000000000000010010000000101110101000000011000000000100000100000000",  -- ROS word 612
   "1000000000000111000000000000000000000000000000010010000000101110101000000001000000000100000000000000",  -- ROS word 613
   "0000001011000000000000000000000000000000000000001110100100000000000000000000000000000000000001000000",  -- ROS word 690
   "0000000000000000000010000000000000000000000000001110100100000000000000000000000000000000000100000000",  -- ROS word 691
   "0000000000000000000010000000000000000000000000010010011000000000000010000000000000000000000100000000",  -- ROS word 692
   "0000000000000000000010000000000000000000000000010010011000000000000010000000000000000000000100000000",  -- ROS word 693
   "1000000000000111100010000000000000000000000000001110001000000100000000000000000000000000000000100000",  -- ROS word 710
   "0000000000000110000000101110010000000000000011001101101000001100000001011100000000000000000000100000",  -- ROS word 711
   "1000000000000000000010000000000000000000000101001110001000000100000010000000000100000100010110100000",  -- ROS word 712
   "1000000000000000000010000101101000000000000000001011101000100000010010000000000000000100000100000000",  -- ROS word 713
   "1000000000000111100010000000000000000000000000001001010110000010000100000000000000000000110000100000",  -- ROS word 790
   "1000000000000111000010101110010000000000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 791
   "1000000000000111100010000000000000000000000000001111000100000100000010000000000000000000110000100000",  -- ROS word 792
   "0000000000000000000010000000000000000000000101101001100110010000000000000000000000000000000100000000",  -- ROS word 793
   "1000000000000111000010110110001000000000000000001111101001001100001111101100000000000100000100000000",  -- ROS word 810
   "1000001001000100100010000000000000000000000001001010000000000000000010000000000000000100000100000000",  -- ROS word 811
   "1000000000000111000010100110000000000000000011001010000100000011000100111100110000000100000100000000",  -- ROS word 812
   "1000001001000100111100000101101000000000000001000111010000000000000010000000100000000100000000000000",  -- ROS word 813
   "1000000000000000000010000000000000000000000000010111000100000001011000000000000000000100000100000000",  -- ROS word 890
   "0000000000000111100010000000000000000000000000000111000000000100000000000000000000111100000000000000",  -- ROS word 891
   "0000000000000000000000000001000000000000000000010001000110000100101010000000000000000100000100000000",  -- ROS word 892
   "1000000000000111100010000000000000000000000000010001001000000100000000000000000000100100010100000000",  -- ROS word 893
   "0000000000000000000010000000000000000000000000010001101000000100101110000000000100000000010110100000",  -- ROS word 910
   "1000000000000000000010000000000000000000000000010001101000000000101110000000000100000100010110100000",  -- ROS word 911
   "1000001010000000000010000010100101110000000000010010000110000100000000000000000000000000000011100000",  -- ROS word 912
   "1000000000000000000010000000000000000000000000000111010000000000000000000000000000000100000100000000",  -- ROS word 913
   "1000000000000000000010000010100000000000000101110010000110000100000000000000000000000100000100000000",  -- ROS word 990
   "0000000000000000000010000101101000000000000011010010101000000100000010000000100000000100000000000000",  -- ROS word 991
   "1000000000000000000010000010100000000000000101110010000110000100000000000000000000000100000100000000",  -- ROS word 992
   "1000000000000000000010000000000000000000000101110010101000000000000010000000000000000100000100000000",  -- ROS word 993
   "1000000000000000001000000000000000000000000000110100001110000100000000000000000000000000000100000000",  -- ROS word a10
   "0000000000000000000000000000000010110000000000010100001010000000000000000000000000000100000100000000",  -- ROS word a11
   "1000000000010000000010000000000000000011010110110100001000000100000010000000000000000100000100000000",  -- ROS word a12
   "0000000000000000000010000000000000000000000010110100001000000001011100000000000000000000000100000000",  -- ROS word a13
   "1000000000000000011110000110010000000000000000010101000110000000000010000000110000000100000100000000",  -- ROS word a90
   "1000000000000111000000011000000000000000000000010101001000000100000010110100001010000110000000000001",  -- ROS word a91
   "0000000000000000000000000100000000000000000000010100100010000100000010000000000000000100000100000000",  -- ROS word a92
   "1000000000000000000000000011010000000001111000010101001010000000000000000000000000000000000100000000",  -- ROS word a93
   "0000000000000000000010000000000000000000000000010110000001000000000010000000000000000000000100000000",  -- ROS word b10
   "0000000000000000000000111000000000000000000000010110000101000001100100000000000000000100000100000000",  -- ROS word b11
   "1000001010000100100010000000000000000000000001010110001010000000000000000000000000010100010100000000",  -- ROS word b12
   "0000000000000010000010000101001000000000000000010110001110000010001000000000000000000100000001000000",  -- ROS word b13
   "1000000000000000000010000110000000000000011000010111001000000000000010000000000000000100000100000000",  -- ROS word b90
   "1000000000000010011110000110110000000011011000010111001000000100000000000000100000011100000111100000",  -- ROS word b91
   "0000000000010010011100000101100000000011010000010111001010100000000010111100110000000110000101000000",  -- ROS word b92
   "0000000001000111000000000110111000000000000000010111001010000000000001001100000000011110110100000000",  -- ROS word b93
   "0000000000010111100001000110101000010101011000011000000110000100000011001000100001000100110100110000",  -- ROS word c10
   "1000000000010111100011000110101000000101011000011000000110000100000011001000100001000100110100110000",  -- ROS word c11
   "1000001011000101000010000110010000000011011000111000100110000000000010000000000000000001011000000000",  -- ROS word c12
   "0000000000000010010111000110011000001101100000011000100111011100000001001010100001000001011100000000",  -- ROS word c13
   "1000001011001100000001111111101010000000000000011001011100000000000011010011101011000000000101100000",  -- ROS word c90
   "1000000001000000000000000001000000100000000101011000101000000100000010000000000000111100000000000000",  -- ROS word c91
   "1000001011001100000010000111101000000000000000011001011100000000000011001100001010000000000001100000",  -- ROS word c92
   "0000000001000000000010000001000000000000000101011000101000000100000010000000000000111100000000000000",  -- ROS word c93
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d10
   "1000000000000010000000000000000000001101001000011010010000100000000000000000000000000000000100110000",  -- ROS word d11
   "0000000000000000000000000000000000000001101000010111011111111100000010000000000000000100000100000000",  -- ROS word d12
   "0000000000010000000010011110010000000100010000011011000010000010001000000000000000000000000100000000",  -- ROS word d13
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d90
   "1000000000000010000010000000000000001100001000011010011000000000000010000000000000000101011111010000",  -- ROS word d91
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d92
   "1000000000010000011110101001111000000101000000011011010100000010001000000000100001000100000100000000",  -- ROS word d93
   "0000000000000000000000000000000000001110000000011011101000000000000000000000000000000100000100000000",  -- ROS word e10
   "1000000000010000000000000110011000000101011000011101001010000000000010000000000000000000000100000000",  -- ROS word e11
   "1000000001000000000000000001001000000000000000111100001110000100000000000000000000110101011000000000",  -- ROS word e12
   "1001010000010010000010000000000000001100110010011100000010000011111010000000000000000000010000000000",  -- ROS word e13
   "1000000000000000000011010000000000000000000000011101001010000100000010000000000000000100000100000000",  -- ROS word e90
   "1000000000001011110110000000000000000000000000011101001000000000000001001100000000000000000000000000",  -- ROS word e91
   "1000000000100111100000000000000000100101010101011100001010000100000010000000000000000000110100110000",  -- ROS word e92
   "1000000000100111100000000001001000100101010101011100001010000100000010000000000000000000110100110000",  -- ROS word e93
   "0011100000000111000010000110110000000000000000011110001010000000000001101100100001000110000000000000",  -- ROS word f10
   "0011100000000111000010000110110000000000000101011110001010000001011011101100100001000110000000000000",  -- ROS word f11
   "1011101011000111000000000110110000000000000001011110001010000100000011101100100001000011101100110000",  -- ROS word f12
   "0011100000000111000010000110110000000000000000111110000010000100000011101100100001000110000000000000",  -- ROS word f13
   "0000000000100000000000000000000000000110011000011110100100000100000010000000000000000100000100000000",  -- ROS word f90
   "0000001011110000000010000000000000000110100000011100010110000010001000000000000000000100000001000000",  -- ROS word f91
   "0000000000100000000000000000000000000110011000011110100100000100000010000000000000000100000100000000",  -- ROS word f92
   "0000000000001011100010000110110000000000000000011111100010000000000001001000100000000010000100000000",  -- ROS word f93
   "1000000000000000000010000000011000000000000000000000011010000100000000000000000000011100000100000000",  -- ROS word 014
   "1000000000000111100010000000000000000000000101000000001010000100000000000000000000000000000011100000",  -- ROS word 015
   "1000000000000100100000000000000000001101101001000000001010000100000010000000000000000000000100000000",  -- ROS word 016
   "1000000000000010000010000010000000001101100000000000001000000000000000000000000000000000000001000000",  -- ROS word 017
   "0000000000000000000000000011010000000000000000001111011100000000000000000000000100000000010110100000",  -- ROS word 094
   "1000000001000000000010000101111000000000000000001001011100000000000010000000000000000100000100000011",  -- ROS word 095
   "1000000000000000000000000011010000000000000000001111011100000000000000000000000100000000010110100000",  -- ROS word 096
   "1000000000000000000000000011010000000000000000001111011100000000000000000000000100000000010110100000",  -- ROS word 097
   "1000000011000000000000000111011000000000000000010010100001111100000000000000000000000100000011100000",  -- ROS word 114
   "0000000001000000000000000000000000000000000000001011001001111100000000000000000000000000000011100000",  -- ROS word 115
   "1000000011000000000000000111011000000000000000010010100001111100000000000000000000000100000011100000",  -- ROS word 116
   "1000000011000000000000000111011000000000000000010010100001111100000000000000000000000100000011100000",  -- ROS word 117
   "1000000000000111000000000110100000010000000000001001001100000000000001001000100000000100000000000000",  -- ROS word 194
   "1000000110000000001000000000011000000000000000001001001000000000000000000000000000000001011111010000",  -- ROS word 195
   "0000000000000111000000000110100000010000000000001001001100000000000001011000100000000100000100000000",  -- ROS word 196
   "1000000000000111000000000110100000010000000000001001001100000000000001010000100000000100000000000000",  -- ROS word 197
   "0000000001100000000001110000000100100010100000000111000101100100000010000000000000000100000100000110",  -- ROS word 214
   "0000000001100000000001111000000100110010100000000111000101100100000010000000000000000100000100000101",  -- ROS word 215
   "1000000001100000000000000000000100000010100000000111000101100100000010000000000000000100000000000100",  -- ROS word 216
   "1000000001100000000001101000000100010010100000000111000101100100000010000000000000000100000000000111",  -- ROS word 217
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 294
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 295
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 296
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 297
   "1000000000000111000010000000000000010000000000010010010100000110001111001000100000000000000000000000",  -- ROS word 314
   "0000000000000000000000111110100000010000000000010001000000000011010110010100100000000000000000000000",  -- ROS word 315
   "0000000000000111000010000000000000010000000000010010010100000110001111011000100000000000000100000000",  -- ROS word 316
   "1000000000000111000010000000000000010000000000010010010100000110001111010000100000000000000000000000",  -- ROS word 317
   "0000001010000010000000000011011000000000000100001011001010000000000010000000000000110000010000000000",  -- ROS word 394
   "1000001010000010000000000011011000000000000100001011001010000000000010000000000000100000010100000000",  -- ROS word 395
   "1000001011010000000000000000000000000011010000000000101010000110100100000000000100000000000101000000",  -- ROS word 396
   "1000001010000010000010000000001000000000000000000101000000000011001110000000000000000001011000000000",  -- ROS word 397
   "0000000000000000000000001000000000000000000101000110001100011001000010000000000000000100000100110000",  -- ROS word 414
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 415
   "0000000000000010000000000111010000000011011000000001101010000100011100000000000000000100000100000000",  -- ROS word 416
   "1000000000000010000010000111010010000011011000000001101010000100011100000000000000000100000100000000",  -- ROS word 417
   "0000000000000010000000000000000000000001111000001001001010000000000010000000000000000000000011010000",  -- ROS word 494
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 495
   "0000000000000010010100000000110000000000000000001011001010000100000000000000100000011100000100000001",  -- ROS word 496
   "1000000000000010000000000111010000000000000000001011001010000100000000000000000000011100000000000001",  -- ROS word 497
   "0000000000000111000000000000000000000000000011001010001010000000000010110100001000000010000000000000",  -- ROS word 514
   "0000000000000010011110000000000000000000000000001010001010000100000010000011111000000100000000000000",  -- ROS word 515
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 516
   "1000000000010111100010000000000000000011010000001010100110100000000000000000000000000100100100100000",  -- ROS word 517
   "1000000000001101000000110000000111100000000000101001000010000000000010000000000000000000000100000000",  -- ROS word 594
   "0000000000000111100010000011011000000000000000010001011100000000000010000000000000000100000011100000",  -- ROS word 595
   "0000000000010000000000000001110000000011010000001000001010000110001110000000000000000100000111010010",  -- ROS word 596
   "0000000000000111100010000100100000000000000000001001001010000100000010000000000000000100000000100000",  -- ROS word 597
   "1000000000000111100010000101011000000011011101001100101010101100000000000000000000000100110100110000",  -- ROS word 614
   "1000000000000000000010000000000000000000000000001100100100101100000010000000000000000100000100000000",  -- ROS word 615
   "1000000000000000011110101000000010000011011000001100010110101100000000000000000000000100000100000000",  -- ROS word 616
   "1000000000000000000010000000000000000000000000001100100100101100000010000000000000000100000100000000",  -- ROS word 617
   "1000000000000111111010000101011000000000000000001101001010000100000010000011100000011000110000110000",  -- ROS word 694
   "1000000000000010011110000000000000000011011000001100010110101100000000000000000000000100100111100000",  -- ROS word 695
   "1000000000000111111000101000000010000000000000001101001010000000000010000011100000011100000000110000",  -- ROS word 696
   "0000000000000010000000000000000000000011011101001100101010101100000000000000000000000100100111100000",  -- ROS word 697
   "1000000000000111000000000110000000000000000000001110001010000000001111110000101000000100000000000000",  -- ROS word 714
   "1000000000000000011000000111000000000000000000001101101010100000000101001111111000000110000000000000",  -- ROS word 715
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 716
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 717
   "0000000000000000000010000000110000000000000000001111001010000000000010000000000000000000000100000000",  -- ROS word 794
   "0000001011000000000010000101111000000000000000001111001010000110101000000000000000000100000001000000",  -- ROS word 795
   "0000000001000000011000000000000000000000000101101101100110000000000000000011000000000000000011100000",  -- ROS word 796
   "1000000001000000011000000000000000000000000101101101100110000000000000000001000000000000000111100000",  -- ROS word 797
   "0000000000000111000010101110100000000000000000010000001011001001001111001100001000000000000100000000",  -- ROS word 814
   "0000001011000000000000000000000000000000000000001100011010000100000010000000001000000000000000000000",  -- ROS word 815
   "1000001011000000000000000000000000000000000000001111101010000000000010000000001000000100000000000000",  -- ROS word 816
   "1000001011000000000000000000000000000000000000001111101010000000000010000000001000000100000000000000",  -- ROS word 817
   "1000000000000111000000110110000000000000000000010001001011001100001111100000001000000100000000000000",  -- ROS word 894
   "1000000000000000000010000000000000000000000100000000101000000100000010000000001000000000000000000000",  -- ROS word 895
   "0000001010000000000010010110111000000000000000000111001010000100000000000000001000000100000000000000",  -- ROS word 896
   "0000001010000000000010010110111000000000000000000111001010000100000000000000001000000100000000000000",  -- ROS word 897
   "1000000000000111000010101110010000000000000011010010001010001100000000000000000000000100000100000000",  -- ROS word 914
   "0000000000000111000010100110000000000000000011010011000000000011000101101000000000000100000000000000",  -- ROS word 915
   "0000000000000000000010000000000000000000000101100000000110010000000010000000000000000000000100000000",  -- ROS word 916
   "1000001010000000000010000010100000000000000000001001001000000000000000000000000000000000000011100000",  -- ROS word 917
   "1000000000000111000000000000000110000000000101110010101010000000000000000001000000000100000000000000",  -- ROS word 994
   "0000000000100000000010000000000110000011010000001110001100101101100100000000000000000000000100000000",  -- ROS word 995
   "1000000000000000000010000000000110000000000101010010101010000100000000000000000000000100000100000000",  -- ROS word 996
   "1000000000000000000010000000000110000000000101010010101010000100000000000000000000000100000100000000",  -- ROS word 997
   "1000000000000000001000000000000000000000000000010100001010000100000000000000000000000000000100000000",  -- ROS word a14
   "1000000000000010000010000000000000010000000000110100001100000000000000000000000010000000000000000000",  -- ROS word a15
   "1000000000000000000010000000000000000000000000010100001010000100000010000000000000000100000100000000",  -- ROS word a16
   "0000000000000000000010000000000000000000000000010100001010000001100010000000000000000000000100000000",  -- ROS word a17
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word a94
   "0000000000000000000010000000000000000000000101010101001010000100000010000000000000000000000100110000",  -- ROS word a95
   "0000000000000000000000000001000000000000000000010000011100000100000010000000000000000100000100000000",  -- ROS word a96
   "0000000000000000000000000011010000000000000011110101001010000000000000000000000100000100010110100000",  -- ROS word a97
   "0000000000010000000010111000000000000011011101010110001010000101100000000000000000000100000001000000",  -- ROS word b14
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b15
   "1000000000000010000010111000000000000000000010010110001101000001100000000000001000000000000000000000",  -- ROS word b16
   "1000001010000000000010000000000000000000000010110101001010000000000000000000000000000000000000001000",  -- ROS word b17
   "1000000001000000000000000011101000000000000001010111001010000000010100000000000000111001011100000000",  -- ROS word b94
   "1000000001100000000010000011110000001011111000010111100010000000000000000000000000011100110100000000",  -- ROS word b95
   "1000000000000010011110000000000000000000000000010111010100000000000010000000100000000000000001100000",  -- ROS word b96
   "0000000000000000000010000111011000000000001000010111001000000100000010000000000000000000000100000000",  -- ROS word b97
   "1000000001000000000011000110110000000000000000011000000100000010001000000000000000000000000001000000",  -- ROS word c14
   "0000000000000111111111000000000000000000000101011000001100000000000011001010100001000010110100110000",  -- ROS word c15
   "0000000000000100100001000101110000000000000000011000000000000011010101001000100101000110000101100000",  -- ROS word c16
   "0000000000000110000010000000000000000000000101011000001010000100000001001100000000000010110100110000",  -- ROS word c17
   "1000000000000010000000000000000000001110010000011001101000010100000000000000000000000001011111010000",  -- ROS word c94
   "0000000001000000000010000001000000000000000000011001001010000000000000000000000000000001011101000000",  -- ROS word c95
   "1000000000000010000000000111101000001101101000011001001100000010001000011100100000000001000101000000",  -- ROS word c96
   "0000000000000010000000000111101000001101101000011001001100000000000011001100100000000101000101000000",  -- ROS word c97
   "1000110000100000000010000000000000000110010000011010010000000100000010000000000000000101000111010000",  -- ROS word d14
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d15
   "1000000000000111000000000111000000001101000000011010001110000000000001001100000000000100000000000000",  -- ROS word d16
   "0000000000000111000010000101101000001101000000011010001101010100000001001100000000000100000000000000",  -- ROS word d17
   "0000000000100000011101010000000000000100000000011010011010100000000010000011100001000100000100000000",  -- ROS word d94
   "1000000000000010000010000000000000001100001000011010011000010100011000000000000000000001011000000000",  -- ROS word d95
   "0000000000000010000010000000000010000000000000011010011010000000000000000000000000000101000000000000",  -- ROS word d96
   "1000000000000010000010000000000000001100001000011010011100000100011000000000000000000010110000000000",  -- ROS word d97
   "1000000000000111100000010000000000000000000000011100000100000010001010000000000000000000110100110000",  -- ROS word e14
   "1011110000000000000010000000000000000000000000011101011100000100000010000000000000011001101001001000",  -- ROS word e15
   "0000000001000000000010000110111000000000000100011100100010000100000010000000000000000100000000001000",  -- ROS word e16
   "1000000000000010000000000000000001011101001000011100001100000000000000000000000000000000010111010000",  -- ROS word e17
   "0000000000000000000010011001111000000000000000011110011100000000000011010000100001000110000000000000",  -- ROS word e94
   "1000000000010000000000000000000000000100111000011111000100000000000010000010100000000000000100000000",  -- ROS word e95
   "1000001001101111000010000101111000000100001000011101000100000011010100000000000000000000000001000000",  -- ROS word e96
   "1010100000100000000000000000000000000100100000011110000010000000000000000000100001000000000100000000",  -- ROS word e97
   "0000000000001011111010011000000000000000000000011110001010000100000000000000000000011000000100000011",  -- ROS word f14
   "1000000000000000011010011000000000000000000000011101011000000000000010000010110000011000000000000011",  -- ROS word f15
   "1010100000000111100010000000000000000000000000011110001100000000000010000000100001000001000000000000",  -- ROS word f16
   "1001010000001010000010000000000000000000000000011110001010000001011010000000000000000100000100000000",  -- ROS word f17
   "0000000000010000011100000010000010000011010000011101010010000000000000000000000000000100000100000000",  -- ROS word f94
   "1000000000000010000010010000000000001110100000011111001100000000000001010000100001000001101001001000",  -- ROS word f95
   "1000001011010111100010000000000000000100100000011111001100000000000010000000000000000101011111010000",  -- ROS word f96
   "0000000001010000000010000000000010000100011000011110100010000100000010000000000000000100000001000000",  -- ROS word f97
   "0000000000000000000000000100110101110000000000001101011010000000101000000000000000000100000100000000",  -- ROS word 018
   "0000000000010000000000000101001000000011010000010100000000000000000000000000000000000100000100000000",  -- ROS word 019
   "0000000000100000001101010000000000000000000000000100000000000011110010000000000000000100000100000000",  -- ROS word 01a
   "1000000000000000000000000100110000000000000000010001010110000100000010000000000000000000000100000000",  -- ROS word 01b
   "0000000000000000011100110000000000000000000000001000000101111101000010000010000000000000000000000000",  -- ROS word 098
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 099
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 09a
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 09b
   "1000000000000000000010000000000000000000000000001011001101111100000000000000000000000100000100000000",  -- ROS word 118
   "0000000001000000000000000000000000000000000000001011001001111100000000000000000000000000000011100000",  -- ROS word 119
   "0000000001000000000000000000000000000000000000001011001001111100000000000000000000000000000011100000",  -- ROS word 11a
   "0000000001000000000000000000000000000000000000001011001001111100000000000000000000000000000011100000",  -- ROS word 11b
   "0000000000000000001000000000000000000001111000001011100110000000000010000000000000000000000011100000",  -- ROS word 198
   "0000000000000010001010000000011000110000000000001001001000000000000000000000000000000001011111010000",  -- ROS word 199
   "0000000000000010001010000000011000110001111000001001001000000000000000000000000000000001011111100000",  -- ROS word 19a
   "0000000000000010001010000000011000110001111000001001001000000000000000000000000000000001011111010000",  -- ROS word 19b
   "0000000000110111100001110000001100100001110101000010000001100111001110000000000000000000000011100110",  -- ROS word 218
   "0000000000110111100001111000001100110001110000000010000001100111001110000000000000000000000011100101",  -- ROS word 219
   "1000000000110111100000000000001100000001110000000010000001100111001110000000000000000000000111100100",  -- ROS word 21a
   "1000000000110111100001101000001100010001110101000010000001100111001110000000000000000000000111100111",  -- ROS word 21b
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 298
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 299
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 29a
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 29b
   "1000000000100000000010001011010000000001110010001000001001111101000010000000000100000100010110100000",  -- ROS word 318
   "0000000000000000000000000011010000000000000010101000001001111100000010000000000100000100010110100000",  -- ROS word 319
   "0000000000000000000000000011010000000000000011101000001001111100000000000000000100000100010110100000",  -- ROS word 31a
   "1000000000000000000000000011010000000000000011101000001001111100000010000000000100000000010110100000",  -- ROS word 31b
   "1000000000000000000010000000000000000000000000000111000010000100000010000000000100000100010110100000",  -- ROS word 398
   "0000001010000000000010000000000000000000000000001000100000000100000010000000000000000100000011100000",  -- ROS word 399
   "0000000000000000000010000000000000000000000000000100010110000000000010000000000100000000010110100000",  -- ROS word 39a
   "0000000000000010000000000000000000000000000000000111001110000100000010000000000000000100010100100000",  -- ROS word 39b
   "0000000000000010000000000000000000000011011000001011001110000000100100000000000000001100000111010000",  -- ROS word 418
   "0000001001000000000010000000000000000000000000101100011100000100000000000000000000000000000100000000",  -- ROS word 419
   "0000000001000000000010000000000001110000000000001110100100000100000010000000000000111001011100000000",  -- ROS word 41a
   "0000001011000000000010000000000001110000000000001110100100000100000010000000000000000000000100000000",  -- ROS word 41b
   "1000000000000111000000000110100000010001111000001001001100000000101110110000100000000100000000000000",  -- ROS word 498
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 499
   "1000001010000000000010000010100000000000000000001001001000000000000000000000000000000000000011100000",  -- ROS word 49a
   "0000000000000000000010000000000000000000000000010011101000000000000011101000000000000100000000000000",  -- ROS word 49b
   "1000000000000000000010000000000000000000000000001100001100001010101000000000000000000100000100000000",  -- ROS word 518
   "1000000000000000000010000000000000000000000000001101001100010000000000000000000000000100000100000000",  -- ROS word 519
   "0000000000000111100010000000000000000000000000001100001100001010101000000000000000000100000000100000",  -- ROS word 51a
   "1000000000000111100010000000000000000000000000001101001100000000000000000000000000000000000000100000",  -- ROS word 51b
   "0000000000000000001000000000000000000000000000001111100000000000000010000000000000000100000100000000",  -- ROS word 598
   "1000000000000111111010000000000000000000000000110001101010001001001111001111110000000010110000100000",  -- ROS word 599
   "0000000000000111100010000000000000000000000101001011011100000100000000000000000000011000000100110000",  -- ROS word 59a
   "1000000000000000000010000100100000000000000000000000001110000000000010000000000000000100000100000000",  -- ROS word 59b
   "1000000000000100100010000000000110000000000000001010100000000000000010000000000000000100000100000000",  -- ROS word 618
   "0000000000000100100010000000000110000000000000001010100100000000000010000000000000000000000100000000",  -- ROS word 619
   "1000000000000100100010000000000110000000000000001001011000000000000000000000000000000100000100000000",  -- ROS word 61a
   "1000000000000100100010000000000110000000000000001010011000000000000000000000000000000100000100000000",  -- ROS word 61b
   "1000000000000100100010000000000110000000000000000000001110000000000010000000000000000100000100000000",  -- ROS word 698
   "1000000000000000000000000101111000000000000000010010000000000011110100000000000000000000000100000000",  -- ROS word 699
   "1000001001000100100010000000000000000000000000010010001100000000000000000000000000000100000100000000",  -- ROS word 69a
   "0000000000100000000010000101101000000011010000001110001100101101100100000000000000000000000100000000",  -- ROS word 69b
   "1000001010000000000010000000000101110000000000001001001000000000000000000000000000000000000011100000",  -- ROS word 718
   "0000001010000000000000000010101101110000000000001001001000000000000000000000000000000000000011100000",  -- ROS word 719
   "1000001010000000000010000010100101110000000011001001001000000000000000000000000000000000000011100000",  -- ROS word 71a
   "1000001010000000000010000010100101110000000000001001001000000000000000000000000000000000000011100000",  -- ROS word 71b
   "0000000000000000000010000000000000000000000000001101001100000000000010000000000000000100100000000000",  -- ROS word 798
   "0000000000100000000010000101101110000011010000001110001100101101100100000000000000000000000100000000",  -- ROS word 799
   "0000000000100000000010000101101000000011010000001110001100101101100100000000000000000000000100000000",  -- ROS word 79a
   "0000000000100000000010000101101000000011010000001110001100101101100100000000000000000000000100000000",  -- ROS word 79b
   "1000001001000000000010000000000000000000000000001010100000000000000010000000000000000100000100000000",  -- ROS word 818
   "0000001001000000000010000000000000000000000000001010100100000000000010000000000000000000000100000000",  -- ROS word 819
   "1000001001000111000000000000000110000000000000000000001110000000000000000000000000000000000100000000",  -- ROS word 81a
   "0000001001000111000000000000000110000000000000001000001110000000000000000000000000000100000100000000",  -- ROS word 81b
   "1000000000000000001000000010010000000000000000001011100110000000000010000000000000000000000100000000",  -- ROS word 898
   "1000000000000000000010000000000000000000000000110000001100010010101000000000000000000100000100000000",  -- ROS word 899
   "0000000001000111000010000000000000000000000000010000100110000000000001001100000000000110000011010000",  -- ROS word 89a
   "1000000000000000000010000000000001100000000000001111001100100010100010000000000000000100000100000000",  -- ROS word 89b
   "1000000000000111000000110110000000000000000011010010001101001100001111110000000000000100000000000000",  -- ROS word 918
   "1000000000000000000010000000000000000000000101110011001100000100000010000000000000000100000100000000",  -- ROS word 919
   "0000000011000000000010000100100000000000000101110001001100000100000010000000000000000000000100000000",  -- ROS word 91a
   "0000000011000000000010000100100000000000000101110001001100000100000010000000000000000000000100000000",  -- ROS word 91b
   "1000000000000000000010000001001000000000000000001101001100100000000010000000000000000000100000000000",  -- ROS word 998
   "1000000011000000000010000000000000000000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 999
   "0000001001000100100010101000000000000000000000001010001110000100000010000000000000000000000100000000",  -- ROS word 99a
   "1000000000000000000010000000000000000000000000001101001110000000000000000000000000000100000100000000",  -- ROS word 99b
   "0000000000000000000010000000000000000000000110110100001100000000000010000000000000111100000000000000",  -- ROS word a18
   "1000001011000000000000000000000000000000000011110100001100000100000000000000000000000100000001011000",  -- ROS word a19
   "1000001011000000000000000000000011000000000000110100001100000100000010000000000000000001000101011000",  -- ROS word a1a
   "0000000000000111100000000000110011010000000000000000000110000000000000000000000000100101000100000000",  -- ROS word a1b
   "0000000000001000000000000000000000000000000000010101001110000000010100000000000000000100000100000000",  -- ROS word a98
   "1000000000001101000010000110010000000000000000110101001100000100000010000000000000000100000100000000",  -- ROS word a99
   "1000000000101000000010000000100000001011110000010111001100000100010100000000000000111000000000000000",  -- ROS word a9a
   "1000000000000111000010000000000010000000000000010101010111010100000010000010100000000100000100000000",  -- ROS word a9b
   "1000000000000111100010000000000000000000000100010110001000000100000000000000000000000100110100110000",  -- ROS word b18
   "1000001010000000000010000000000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word b19
   "0000000000000111100010000000000000000000000000010110001010000000000000000000000000000000110100110000",  -- ROS word b1a
   "0000000000000111000000000110110000000000000000010111011100000100000000111100110000000100000100000000",  -- ROS word b1b
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b98
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b99
   "0000000000000000000010000000000000000000000000010111001100000100000000000000000000000000000100000000",  -- ROS word b9a
   "1000000000000010011110000000000000000000000000010111001110000000000000000000100000000000000000000000",  -- ROS word b9b
   "0000000000000110011111000110110000000000000000011000001110000000010011110110100001000000000100001000",  -- ROS word c18
   "1000000000000000000000100000000000000000000000111000001100000100000010010110100001000010000100000000",  -- ROS word c19
   "0000000000000110011111000110110000000000000101111000001110000000010011110110100001000100110000110000",  -- ROS word c1a
   "0000001001100000010100010110111000000010001000011000011010000000000000000010000000000000000000000000",  -- ROS word c1b
   "1000000000101111010110000110110000000011010000011001001110000100000001001100100000000010000000000011",  -- ROS word c98
   "0000000000101111010110000110110000000011010000011001001111000110001001001100100000000110000000000011",  -- ROS word c99
   "0000000001000000000010000110111000000000000000010111011101111100000000000000000000000100000000000010",  -- ROS word c9a
   "0000000001110000000010000110001000001000010000010111010101111100000000000000000000000000000100110000",  -- ROS word c9b
   "0000000000010000000000000000000010000011010000011010001100000000000010000000000000000100000100000000",  -- ROS word d18
   "1000001010000000000010000000000000000000000000011010001000000000000010000000000000000000000001000000",  -- ROS word d19
   "1000001010000000000010000000000000000000000000011010001000000000000010000000000000000000000001000000",  -- ROS word d1a
   "1000001010000000000010000000000000000000000000011010001000000000000010000000000000000000000001000000",  -- ROS word d1b
   "0001010000001011111100000101011000000000000000011011001100000100000000000000100000000000000001001000",  -- ROS word d98
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d99
   "1000001011001101000010000000000000000000000000111011001110000001001100000000000000000000000011010000",  -- ROS word d9a
   "1000000000000010000010000111011000001100011000011010000010000000010101001100100000000100000100110000",  -- ROS word d9b
   "1000000000010010000010000110011000000101011000011101011111010100000000000000000000000000010000000000",  -- ROS word e18
   "1000000000010000000010000001000000000100111000011100011010000110001010000010100000000100000100000000",  -- ROS word e19
   "1000000001000000000000000000101000000000000100011100001100000100000010000000000000000100000000001000",  -- ROS word e1a
   "1000001010000000000010000000000000001100101000111100000100000100010101001000100000000100000101000000",  -- ROS word e1b
   "1000000000010010000010000101111000000011010000010101011010000100000000000000000000000001101001001000",  -- ROS word e98
   "1000000000000010011100000000000000001100010000011100011100000010001000000000000000000100010000000000",  -- ROS word e99
   "0000000000000011100000000000000000001100101000111100010100000100000010000000000000000100110100110000",  -- ROS word e9a
   "0000001011001111010101000101101011010000000000011101010111010100000010000010100001110000000000000000",  -- ROS word e9b
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word f18
   "0000000000001111000011010101101000000000000000011110000100100010001000000000000000000100000000001011",  -- ROS word f19
   "0000000000000110000010000110110000000000000011011110001100000100000010000000000000000100000001000000",  -- ROS word f1a
   "0000000000000111000000000000000000000000000011011110001110000010001010000000000000000100000100000000",  -- ROS word f1b
   "0000000000000010000000001000000000001100111000011111001110000010001001010000100001000100000100110000",  -- ROS word f98
   "0000000000000010000000000000000000001100000000011111010000000011111010000000000000000100000100000000",  -- ROS word f99
   "1000000000000010000010000000000000001100111000011111001110000000000000000011110000000100000100110000",  -- ROS word f9a
   "1000001011000111100000000000000000000000000000011000010010000100000000000000000000000001000111010000",  -- ROS word f9b
   "0000000000000000000000110110001001100000000000000000001111001100001111110000000000000000000000000000",  -- ROS word 01c
   "0000001010000000000010000000000000000000000100010001001100000000000010000000000000110100010000000000",  -- ROS word 01d
   "1000000000000000000010000000000000000000000000010011001100000000000100000000000000000100000100000000",  -- ROS word 01e
   "1000000000000000000010000000000000000000000000010011001100000000000100000000000000000100000100000000",  -- ROS word 01f
   "0000000001110000000010000110001000001000010000010111010101111100000000000000000000000000000100110000",  -- ROS word 09c
   "0000000001110000000010000110001000001000010000010111010101111100000000000000000000000000000100110000",  -- ROS word 09d
   "0000000001110000000010000110001000001000010000010111010101111100000000000000000000000000000100110000",  -- ROS word 09e
   "0000000001110000000010000110001000001000010000010111010101111100000000000000000000000000000100110000",  -- ROS word 09f
   "0000000000010000000001000110111000000001100000001011001011111100000000000000000000000100000100000000",  -- ROS word 11c
   "1000000110100000000001000000010000000001100000001000001101111100000000000000000000000100000011010000",  -- ROS word 11d
   "0000000001000000000000000000000000000000000000001011001001111100000000000000000000000000000011100000",  -- ROS word 11e
   "0000000001000000000000000000000000000000000000001011001001111100000000000000000000000000000011100000",  -- ROS word 11f
   "0000000000100000000001000110111000000001100000001001000011111100000000000000000000000100000100000000",  -- ROS word 19c
   "1000000000000000000010000000000000000000000000001000000001111100000000000000000000000100000100000000",  -- ROS word 19d
   "0000000110000010001010000000011000000001111000001001001000000000000000000000000000000001011111100000",  -- ROS word 19e
   "0000000110000010001010000000011000000001111000001001001000000000000000000000000000000001011111010000",  -- ROS word 19f
   "1000000000110111100001110000001100100001110101000010000001100111001110000000000000000000000100000110",  -- ROS word 21c
   "1000000000110111100001111000001100110001110000000010000001100111001110000000000000000000000100000101",  -- ROS word 21d
   "0000000000110111100000000000001100000001110000000010000001100111001110000000000000000000000000000100",  -- ROS word 21e
   "0000000000110111100001101000001100010001110101000010000001100111001110000000000000000000000000000111",  -- ROS word 21f
   "1000001001000100100000000101111000000000000000000100000110000100000010000000000000000000000100000000",  -- ROS word 29c
   "1000001001000100100000000101111000000000000000000100000110000100000010000000000000000000000100000000",  -- ROS word 29d
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 29e
   "0000000000000100100000000101111000000000000100000111011010000100000000000000000100000100010110100000",  -- ROS word 29f
   "1000000001010000000000000111000011010011010000010001010100000000000000000000000000000100000001000000",  -- ROS word 31c
   "0000000000000111000000000000000000000000000000010001001110000000000001001100000000000000000000000000",  -- ROS word 31d
   "0000000000000000000010000111100000000000000000001011000010100000000000000000000000000000000100000000",  -- ROS word 31e
   "0000000000000000000010000111100000000000000000001011000010100000000000000000000000000000000100000000",  -- ROS word 31f
   "1000001010000010000010000000001000000000000000000101000000000011001110000000000000000000000001000110",  -- ROS word 39c
   "1000000000110111100010000000001000000001110101000010000000000011001110000000000000000101011111100000",  -- ROS word 39d
   "0000001010000010000010000000001000000000000000000101000000000011001110000000000000000000000100000110",  -- ROS word 39e
   "0000000000000000000010000000000000000000000000010011010110000000011100000000000000000000000111010001",  -- ROS word 39f
   "0000000000000000000000110110001001100000000000001000001111001100001111100000000000000100000100000000",  -- ROS word 41c
   "0000001010000000000010000000000000000000000100010001001100000000000010000000000000110100010000000000",  -- ROS word 41d
   "1000000011000000000010000000000000000000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 41e
   "1000000011000000000010000000000000000000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 41f
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 49c
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 49d
   "0000000000000000000000000001001101100000000000001101001100100000000010000000000000000000100000000000",  -- ROS word 49e
   "0000000011000000000000000000000101100000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 49f
   "0000000000000010001000000000000000000001101000001001001000000000000000000000000000000001011000000000",  -- ROS word 51c
   "1000001101000010000010000000011000000001111000001000011110000000000000000000000100001000000011100000",  -- ROS word 51d
   "1000000000000111100010000000000000000000000000010011001010010101100100000000000000000100110100110000",  -- ROS word 51e
   "1000000000000111000000000000000000000000000000001011010100000000100100000000000000000000000100000000",  -- ROS word 51f
   "0000001011011101000010000001001000000011010000001000001100000100001000000000000000000000000100000000",  -- ROS word 59c
   "0000000001011101000000000000000000000001100000001000001100000100000010000000000000000000000001000000",  -- ROS word 59d
   "0000001001000010000000000000000000000000000000001010010001001000000000000000000000000001011000000000",  -- ROS word 59e
   "0000000000000010000000000000000000000000000000001111100100000000000010000000000000000001011000000000",  -- ROS word 59f
   "1000000000000010000010000111011000000000000000001100010000000000000010000000000000000100000100000000",  -- ROS word 61c
   "0000000000000111000010000110010000000000000000001100001000000000000001001100000000000010000100000000",  -- ROS word 61d
   "0000000000000111100010000000000000000000000000001111011000000000001110000000000000011000000100110000",  -- ROS word 61e
   "0000000000100000000010000111111000000011010000010001011000000000000010000000000000000000000100000000",  -- ROS word 61f
   "1000000000000111100010000000000000000000000000001101001110000000000010000000000000000000110000100000",  -- ROS word 69c
   "0000000000000111100010000000000000000000000101001101001110000100000010000000000000000100000000100000",  -- ROS word 69d
   "1000000000000111100010000000000000000000000000001010001100000101001110000000000000000000110000100000",  -- ROS word 69e
   "0000000000000000011010000000000000000000000000001010001100000001001111101111110000000110000000000000",  -- ROS word 69f
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 71c
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 71d
   "0000000000000000000000000001001101100000000000001101001100100000000010000000000000000000100000000000",  -- ROS word 71e
   "0000000000000000000000000000000101100000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 71f
   "0000001001000000000010000000000110000000000000001000000000000011001100000000000000000000000100000000",  -- ROS word 79c
   "0000000001000000000000000000000110000000000000000110000000000011001110000000000000000000000011100000",  -- ROS word 79d
   "0000001011000000000000000000000000000000000000001111001110000000010010000000000000000000000001000000",  -- ROS word 79e
   "0000000000000000000010000000000000000000000000001111001110000000000000000000000000000000000100000000",  -- ROS word 79f
   "0000000000000111100010000000000000000000000101001011011100000100000000000000000000000000110100110000",  -- ROS word 81c
   "0000000000100000000010000111111000000011010000010001011000000000000010000000000000000000000100000000",  -- ROS word 81d
   "1000000000000000000000000101100011000000000000001110000010000100000000000000000000000000000100000000",  -- ROS word 81e
   "1000000000000000000000000001000011000000000110100100101000000000000010000000000000000000000100000000",  -- ROS word 81f
   "1000000000000000000010000101011000000000000000010010001110000011000110000000000000000000010000000000",  -- ROS word 89c
   "1000001010000000000010000101101000000000000000010001001110000100000000000000000000000100010111010000",  -- ROS word 89d
   "1000000000000000000000000110001101110000000101010001001110000100000010000000000000000000000100000000",  -- ROS word 89e
   "0000000000000000000010000000000000000000000000001111001110000100000010000000000000000000000100000000",  -- ROS word 89f
   "0000001010000101000000000111011110000000000000001011010001000000000010000000000000000100010111010000",  -- ROS word 91c
   "0000001010000101000000000111011110000000000000001011010001000000000010000000000000000100010111010000",  -- ROS word 91d
   "0000001010000100000000000000000110000000000000001011010001000000000010000000000000000100010111010000",  -- ROS word 91e
   "0000001010000100000000000000000110000000000000001011010001000000000010000000000000000100010111010000",  -- ROS word 91f
   "1000000000100000000000000110110000000001100000010011001110000000000010000000000000000000000100000000",  -- ROS word 99c
   "0000000000000011000000001000000000000000000000010011001110000100000000000000100000000000000000110000",  -- ROS word 99d
   "1000000000000000000010001110111000000001111000010011001110000100000010000000000000000100000100000000",  -- ROS word 99e
   "1000000000100000000000000111011000000001110000001111100100000100000000000000000000000000000100000000",  -- ROS word 99f
   "1000000000010010000010000000000000010011010000110100001110000000000010000000000010000000000000000000",  -- ROS word a1c
   "0000000000000000000010000000000000000000000110110100000010000100000000000000000000000000000100000000",  -- ROS word a1d
   "1000000000000010000010000000000001000011011000110100001000000100000000000000000010000000000000000000",  -- ROS word a1e
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word a1f
   "1000000000000000000010000100010000000000000000010101001000000000000000000000000000000100000100000000",  -- ROS word a9c
   "0000000000000000000000000100000000000000000000010101001000000000000000000000000000000100000100000000",  -- ROS word a9d
   "0000000000000000011101110000000000000011111000010101100000000100000010000000100001000100000100000000",  -- ROS word a9e
   "1000000000000000011110000011010000000000000000010101010000000000000010000010000000000000000000000000",  -- ROS word a9f
   "0000000000000000000000000000000011010000000000010100010000000000000010000000000000000100000100000000",  -- ROS word b1c
   "1000000000001001100010000000001000000000000000010110010110000000000000000000000000000100000100000000",  -- ROS word b1d
   "1000001001000000000000000000000010110000000000110110001110000100000010000000000000000000000100000000",  -- ROS word b1e
   "0000000000000010000010000000000001000011011001010110010110000100000000000000000010000100000000000000",  -- ROS word b1f
   "1000000000000111000000000000000000000000000000010111001110000000000011101100000000000110000000000000",  -- ROS word b9c
   "0000000000000000000010000000101000000000011000010111001110000100000010000000000000000000000100000000",  -- ROS word b9d
   "1000000000000000000010011000000000000000000000010111100110000000000000000000001010000000000000000001",  -- ROS word b9e
   "0000000000000000000000000011101000000000001001010111010000000000000000000000000000000100000100000000",  -- ROS word b9f
   "1000000000010000011011001000010000000101011000011000000100000100000000000011100001000100000100000000",  -- ROS word c1c
   "1000000001110000010100000110011000000101000000011000011100000000000010000000000000000100110000001000",  -- ROS word c1d
   "0000000000000000010101000110011000000000000000011000000010000110001001001010100000000100000100000000",  -- ROS word c1e
   "0000000001100000000000000100011000000101000000011001000000000100000000000000000000000100000100110000",  -- ROS word c1f
   "0000000001010000000010000110011000010101010000011000011000001110100010000010110000111000000100000000",  -- ROS word c9c
   "0000000001010000000010000110011000010101010000011000011000001110100010000010110000111000000100000000",  -- ROS word c9d
   "0000000001000000011000000110110000000000000000011001010000000110000101110100110100000010000011100000",  -- ROS word c9e
   "0000000001010000000010000110011000010101010000011000011000001110100010000010110000111000000100000000",  -- ROS word c9f
   "1000001001010010000000000110011000000101010000011011101010000100000010000000000000000000000100000000",  -- ROS word d1c
   "1000000000010000000010000101101000000011010000011010001101010100010100000000000000000100000100000000",  -- ROS word d1d
   "0000000000000000000000000001111000001100100000011010001110000010001010000000000000000000000001000000",  -- ROS word d1e
   "1000000000000111000000000000000000000000000010011010010110000000000001001100000000000000000100111000",  -- ROS word d1f
   "0000000000001100000000000110100000001101001000011011001110000100000000011100000000000110000110001000",  -- ROS word d9c
   "1000000000001100000000000110100000001101001000011011001110000100000000011100000000000110000010011000",  -- ROS word d9d
   "1000000000000110000010000110011000000000000000011011001110000100000011001110110000000001011000000000",  -- ROS word d9e
   "1000000001000111000010000110110000000000000000011011010000000000000000000010110000000001000011100000",  -- ROS word d9f
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word e1c
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word e1d
   "0001010001000000000000110000000000000000000000011100010000000011111010000000000000000101011101000000",  -- ROS word e1e
   "0000000000010000000010000000000000000100110100011101011000000100000010000000000000000000000100000000",  -- ROS word e1f
   "0000000000000000000010011101101000000000000111011101000010000000000010000000000000000000000100000000",  -- ROS word e9c
   "1000000000000000000010011101101000000000000111011101000010000000000010000000000000000001101000000000",  -- ROS word e9d
   "0000000000100000000000000000000010000100101000011101010010000100000010000000000000000100000100000000",  -- ROS word e9e
   "1000000000000010000000000000000000001100110000011101001110000100000000000000000000000100000001000000",  -- ROS word e9f
   "1010100000001111000010000110110000000000000000011110001110000100101110000000100001000100000100000000",  -- ROS word f1c
   "1000000000000000010100100110011000000000000101011101010100000000000010000000100001000000000100000000",  -- ROS word f1d
   "0000000000000111100011010101101000000000000000011110000100100010001000000000000000000101101000110000",  -- ROS word f1e
   "1000000000000000000011010000000000000000000101011110010000000000000000000000000000000001101000110000",  -- ROS word f1f
   "0000000000000010000000011110101000001110001000011111001110000110001001010000100001000001011000000000",  -- ROS word f9c
   "1010100000001111000010000110101000000000000000011110100100000000000010000000100001000000000000001011",  -- ROS word f9d
   "0010101101000000000000000000000000000000000000011110101000000010001001010000100001000100000100000000",  -- ROS word f9e
   "1010100000001111000010000001001000000000000000011110100100000000000010000000100001000000000000001011",  -- ROS word f9f
   "1000000000000000000010000000000011110000000000010000000100000011001100000000000000000100000100000000",  -- ROS word 020
   "1000000000000111111010000000000000000000000000110001101010001001001111001111110000000010110000100000",  -- ROS word 021
   "0000000000000000000000000000001000000000000101000010000000000011001110000000000000000100000100110000",  -- ROS word 022
   "1000000000000111000000000100100000000000000000101000001110000000000000000000000000000000000100000000",  -- ROS word 023
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a0
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a1
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a2
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a3
   "1000000000100000000000000011010000000001000010010011010011111100000000000000000100000000010110100000",  -- ROS word 120
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 121
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 122
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 123
   "1000001011010000000010000000010000000010000000000100100011111100000010000000000000000000000011100000",  -- ROS word 1a0
   "1000001011010000000010000000010000000010000000000100100011111100000010000000000000000000000011100000",  -- ROS word 1a1
   "1000001011010000000010000000010000000010000000000100100011111100000010000000000000000000000011100000",  -- ROS word 1a2
   "1000001011010000000010000000010000000010000000000100100011111100000010000000000000000000000011100000",  -- ROS word 1a3
   "1000000011110111111111110000001100100001110101000001000001100111001110000011110000000000000011100110",  -- ROS word 220
   "1000000011110111111111111000001100110001110000000001000001100111001110000011110000000000000011100101",  -- ROS word 221
   "0000000011110111111110000000001100000001110000000001000001100111001110000011110000000000000111100100",  -- ROS word 222
   "0000000011110111111111101000001100010001110101000001000001100111001110000011110000000000000111100111",  -- ROS word 223
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a0
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a1
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a2
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a3
   "1000000000000010011010000000000011100000000000000111000000000100000010000000000010000000000000000000",  -- ROS word 320
   "0000000000000010011010000000000011100000000000000111011010000100000010000000000010000100000000000000",  -- ROS word 321
   "1000000000000010011010000000000011100000000000000111100110000000000010000000000010000000000000000000",  -- ROS word 322
   "1000000000000000000000000000000011100000000000000110010110000000000000000000000000000000000100000000",  -- ROS word 323
   "1000000000000000000010000000000000000000000101010000001000100000000010000000000000000100000100000000",  -- ROS word 3a0
   "1000000000000111000000000000000000000000000000001110101000000000000001001100000000000010000100000000",  -- ROS word 3a1
   "0000000000000000000000000000000110010000000101000110011000000000000000000000000000000100000100000000",  -- ROS word 3a2
   "1000000000000000000010000000000010100000000000010101001110000100000010000000000000000100000100000000",  -- ROS word 3a3
   "0000000000000010000010000110101010000000000000000110001110000000000010000000000000000100000001000000",  -- ROS word 420
   "0000000000000010000010000110101010000000000000000110001110000000000010000000000000000100000001000000",  -- ROS word 421
   "0000000000000010000010111110101000000000000000001001010001000010001000000000000000000100000001000000",  -- ROS word 422
   "1000000000000010000000111110101011010000000000001001010001000010001000000000000000000100000001000000",  -- ROS word 423
   "1000000000000000000010011101101000000000000000010011001110000000000000000000000000000100000100000000",  -- ROS word 4a0
   "1000000000000110000010000000000001010000000000010001001110000010000101001100000000011000000000110000",  -- ROS word 4a1
   "1000000000000000000010011000000000000000000000010011001110000000000000000000000000000100000100000000",  -- ROS word 4a2
   "0000000000000000000010000000000000000000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 4a3
   "0000000000000110000000111110110000000000000011001000000110000000000001001100000000011000000000110000",  -- ROS word 520
   "1000000000000000000010000110110000000000000011001011001100000100000000000000000000000100000100000000",  -- ROS word 521
   "0000000000000111000010111000000000000000000101101010010001000000000011001100000000000100000000000000",  -- ROS word 522
   "0000000000000000000010000000000000000000000011010010011000000000000010000000000000000000000100000000",  -- ROS word 523
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 5a0
   "1000001010000000011100000110111101100000000100101000010000100000001110000000100000000100010001000000",  -- ROS word 5a1
   "1000000000000111000000000101110000000000000000001011010000000000000010000000000000000000000100110000",  -- ROS word 5a2
   "1000000000000000011110000110111000000000000000001000010000000100000000000000100000000000000000000000",  -- ROS word 5a3
   "1000000000000010000010000111011000000000000000001100010000000000000010000000000000000100000100000000",  -- ROS word 620
   "0000001011000111000010000000000000000000000000001100010000000100000001001100000000000110010000000000",  -- ROS word 621
   "1000001010000000000010000000000101110000000100001100010000000100000010000000000000000100010111100000",  -- ROS word 622
   "0000000000000000000000000001110000000000000000000111011100000000000000000000000100000100010110100000",  -- ROS word 623
   "1000000000000000000010011000000000000000000000000001101000000000000010000000000000000100000100000000",  -- ROS word 6a0
   "1000000000000000000010011110001011010000000000000001101000000000000010000000000000000100000100000000",  -- ROS word 6a1
   "1000000000000000000010011110001011010000000000000001101000000000000010000000000000000100000100000000",  -- ROS word 6a2
   "1000000000000000000010011000000000000000000000000001101000000000000010000000000000000100000100000000",  -- ROS word 6a3
   "0000000000000000000010000000000001010000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 720
   "0000000000000000000010000000000000000000000000001100010100100001100000000000000000000000000100000000",  -- ROS word 721
   "1000000000000000000000000000000011010000000000010000001110000000000010000000000000000000000100000000",  -- ROS word 722
   "0000000000000000000010000000000000000000000000001100010100100001100000000000000000000000000100000000",  -- ROS word 723
   "1000000000000111000010000000000000010000000000010010010100000110001110110000100000000000000000000000",  -- ROS word 7a0
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 7a1
   "0000000000000000000010000000000000000000000101101010010100000100000010000000000000000000000100000000",  -- ROS word 7a2
   "0100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",  -- ROS word 7a3
   "0000000000000111000010111110100000010000000011010000010001001001001110110000100000000100000000000000",  -- ROS word 820
   "1000001010000000000000000110010000000000000100001111000100000100000000000000000000010000010100000000",  -- ROS word 821
   "0000000000000000000010000000000000000000000101101010010100000100000010000000000000000000000100000000",  -- ROS word 822
   "0000000000000000000010000001001000000000000101101010010100000100000010000000000000000000000100000000",  -- ROS word 823
   "1000000000000111000000000000000000000000000000001000010110000110001111000100110000000000000100000000",  -- ROS word 8a0
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 8a1
   "0000000000000000000010000000000000000000000101110011010100000101100000000000000000000000000100000000",  -- ROS word 8a2
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 8a3
   "1000000000000111000000111110100000000000000011010010010001001001001111000100110000000000000100000000",  -- ROS word 920
   "1000001010000000000000000110010000000000000100001111000100000100000000000000000000010000010100000000",  -- ROS word 921
   "0000000000000000000010000000000000000000000101110011010100000101100000000000000000000000000100000000",  -- ROS word 922
   "0000000000000000000010000001001000000000000101110011010100000101100000000000000000000000000100000000",  -- ROS word 923
   "0000000000000111000000000000000000000000000000001001010110000110001111101110100000000100000100000000",  -- ROS word 9a0
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9a1
   "0000000000000000000010000000000000000000000101110011010100000101100000000000000000000000000100000000",  -- ROS word 9a2
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9a3
   "1000000000000010000000000000000000000000000000010100010000000110001001001000100000000100000001100000",  -- ROS word a20
   "1000000000000000000000000010000000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word a21
   "1000000000000010000000000000000000000000000000010100010010000010001001001000100000000100000001100000",  -- ROS word a22
   "0000000001100000000010000110010000000001110000010100011000000000000000000000000000011100110011100000",  -- ROS word a23
   "1000000000000000011110010011100010110000000000110101010010000000000000000011100001000100000100000000",  -- ROS word aa0
   "1000000000000000011100000000000000000000000000110101010001000100110111001111110000000010000100000000",  -- ROS word aa1
   "1000000000000000011110010011100010110000000000110101010010000000000000000011100001000100000100000000",  -- ROS word aa2
   "1000000000001000000000000011100010110000000000010101001010010100000000000000000000000000000100000000",  -- ROS word aa3
   "1000000000000000000000111000000000000000000011110110001101000001100000000000000000000000000100000000",  -- ROS word b20
   "1000000000000000000000111000000000000000000011110110010010000101100000000000000000000000000100000000",  -- ROS word b21
   "0000000000000111000000000011101000000000000000010111100100000100000011001111110000000110000100000000",  -- ROS word b22
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b23
   "1000000000000000000010000000000000000000000000010111010000000001101000000000000000000100000100000000",  -- ROS word ba0
   "0000000000000000000010000011110000000000000000010100100010000100000000000000000000000000000100000000",  -- ROS word ba1
   "1000001011000000011110000110101000000000000000010111010000000100000010000000100000000000000001100000",  -- ROS word ba2
   "1000000000000111000000000000000000000000000000010111010010000000000000111100000000000110000000000000",  -- ROS word ba3
   "1000000000010000000000000110011000100101010000011000011000001110100010000000000000000000000100000000",  -- ROS word c20
   "1000110000101111011000010001000000000010001000011000010010111100000011001111110000000011000111010000",  -- ROS word c21
   "0000110000101111011010010000000000000010001000011000010010111100000011001111110000000011000111010000",  -- ROS word c22
   "1000000000010000000000000110011000100101010000011000011000001110100010000000000000000000000100000000",  -- ROS word c23
   "0000000000110000000010000000000000001000010000010101001011111100000010000000000000000000000100000000",  -- ROS word ca0
   "1000000000000000000000000110010000000000000000010101001101111100000010000000000000000000000100000000",  -- ROS word ca1
   "0000000001100000010111000110100000000101101000011001011000000100000001001000100001000100000011100000",  -- ROS word ca2
   "1000000001100000010101100110100000000101101000011001011000000100000001001000100001000100000011100000",  -- ROS word ca3
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word d20
   "0000100001100000000010000000000000000110001000011010001010000000000000000000000000000001000111010000",  -- ROS word d21
   "1000000000001111000010000101101000000000000000011001011110000000000010000000000000011100000100000000",  -- ROS word d22
   "0000100000100000000010000110011000000110011000011010010010000000011000000000000000000001000111010000",  -- ROS word d23
   "1000001010000111000000000000000000000000000000011011010010000011111010000010110000000100010001011000",  -- ROS word da0
   "0000000000000000011100000101011000000000000000011011001100000100000000000000100000000000000001001000",  -- ROS word da1
   "1000001010000000011100110000000000000000000001011011011100000000000000000000100001000100010001001000",  -- ROS word da2
   "1000000000000000000000000111011000001100011011111011011000000000000000000000000000000000000100000000",  -- ROS word da3
   "1000001010000000000010000010111000001100110000011100010000000100000010000000000000000100010101000000",  -- ROS word e20
   "1000001010000000000010000010111000001100110000011100010000000100000010000000000000000100010101000000",  -- ROS word e21
   "1000001010000000000010000010111000001100110000011100001110000100000010000000000000000100010101000000",  -- ROS word e22
   "1000000000010000000010000000000000000100110100111100010010000010001010000000000000000100000100101000",  -- ROS word e23
   "0000000000000000000000011000000010000000000000011101010000100000000000000000000000000100000101001011",  -- ROS word ea0
   "0000000001000000000000000000000000000000000000011101001000000100000000000000000000000100000100110000",  -- ROS word ea1
   "0000000000000010000000000000000000000000000000011101010011010100000010000000000000000100000100110000",  -- ROS word ea2
   "0001011010110000000000000000000000000100110000011100000010000011111010000000000000000100010111010000",  -- ROS word ea3
   "1010100000000000000010000000000000000000000000011110010000000101011010000000100001000100000100000000",  -- ROS word f20
   "1000000000000000000010011000000000000000000011111101011100000000000000000000000000000100000100000000",  -- ROS word f21
   "0000000000000111100010000101101000000000000000011110000100100010001000000000000000000101101000110000",  -- ROS word f22
   "0000000000100111100000000000000000000101011101011110010000000000000010000000000000000100110100110000",  -- ROS word f23
   "0000000000000010000010000000000000001100100000011001101000010100000000000000000000000001011101000000",  -- ROS word fa0
   "1000000000100000000000000000000000000100001000011111001100000100000010000000000000000000000100000000",  -- ROS word fa1
   "0000000000000111100010000000000000000000000000011000010100000000000000000000000000000100000000100000",  -- ROS word fa2
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fa3
   "0000000000000000000000000000001000000000000101000001000000000011001110000000000000000100000100110000",  -- ROS word 024
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 025
   "1000000000000000011110000000111000000000000000010000011100000100000000000010110000000000000000000000",  -- ROS word 026
   "1000000011000000000010000000000001100000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 027
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a4
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a5
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a6
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a7
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 124
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 125
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 126
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 127
   "0000000000100111100010000110011000000010000000010011101011111100000010000000000000000100000011100000",  -- ROS word 1a4
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 1a5
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 1a6
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 1a7
   "0000000011110111111111110000001100100001110101000001000001100111001110000011110000000000000100000110",  -- ROS word 224
   "0000000011110111111111111000001100110001110000000001000001100111001110000011110000000000000100000101",  -- ROS word 225
   "1000000011110111111110000000001100000001110000000001000001100111001110000011110000000000000000000100",  -- ROS word 226
   "1000000011110111111111101000001100010001110101000001000001100111001110000011110000000000000000000111",  -- ROS word 227
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a4
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a5
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a6
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a7
   "0000000000000000000010000000000000000000000000000110010110000000000000000000000000000000000100000000",  -- ROS word 324
   "1000000000000000001000000000000000000000000000100110010110000000000010000000000000000000000100011000",  -- ROS word 325
   "1000000000001011101000011000000000000000000000100110010110000000000010000000000000000000000100000000",  -- ROS word 326
   "1000001010000000001000000000000000000000000000100110010110000000000010000000000000000000000100000000",  -- ROS word 327
   "1000000000000010010110000000000000010000000000100011101000000100000010000000000010000000000000000000",  -- ROS word 3a4
   "0000000000100000010110000000000000000011010000100011101000000100000010000000000000000000000100000000",  -- ROS word 3a5
   "1000000000000010000000000000000000000011011000000111001010000100000010000000000000010000010100000000",  -- ROS word 3a6
   "0000000000000010000000000000000000000011011000000111001010000100000010000000000000000000010000000000",  -- ROS word 3a7
   "1000000000000111000000111110100000000000000011001000010011001001001111101110100000000000000100000000",  -- ROS word 424
   "1000001010000000000000000110010000000000000100001111000100000100000000000000000000010000010100000000",  -- ROS word 425
   "0000000000000000000010000000000000000000000101110011010100000101100000000000000000000000000100000000",  -- ROS word 426
   "0000000000000000000010000001001000000000000101110011010100000101100000000000000000000000000100000000",  -- ROS word 427
   "0000000000000111000000000000000000000000000000001011010110000110001111001100000000000000000000000000",  -- ROS word 4a4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4a5
   "0000000000000000000010000000000000000000000101101000011010000000000000000000000000000000000100000000",  -- ROS word 4a6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4a7
   "1000000000000111000000111110100000000000000011001010010011001001001111001100000000000100000000000000",  -- ROS word 524
   "1000001010000000000000000110010000000000000100001111000100000100000000000000000000010000010100000000",  -- ROS word 525
   "0000000000000000000010000000000000000000000101101000011010000000000000000000000000000000000100000000",  -- ROS word 526
   "1000000000000000000010000000000000000000000101101000011010000000000010000000000000000100000100000000",  -- ROS word 527
   "1000000101000000011100110000000111100000000000000010100100000000000001001110000100000010101100000000",  -- ROS word 5a4
   "1000000101000000011100110000000111100000000000000010100100000000000001001110000100000010101100000000",  -- ROS word 5a5
   "1000000000000000000001000000000000000000000000000011100010000000000010000000000000000000000100000000",  -- ROS word 5a6
   "1000000000000000000001000000000000000000000000000011100010000000000010000000000000000000000100000000",  -- ROS word 5a7
   "0000001001001010000010000110101010010000000000001100011000000000000010000000000000000000000100000000",  -- ROS word 624
   "0000001001001010000011111000000000000000000000010000011110000000000000000000000000000000000100000000",  -- ROS word 625
   "0000000000001010000000000011010010010000000000001111011110000000000000000000000000000100000100000000",  -- ROS word 626
   "0000001001001010000011111000000000000000000000010000011110000000000000000000000000000000000100000000",  -- ROS word 627
   "0000001010001010000000000100110010010000000110000000001100000100011110010000000000000000110000110000",  -- ROS word 6a4
   "1000000000100000000111010000000101110000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 6a5
   "0000001010001010000000000100110010010000000110000000001100000100011110010000000000000000110000110000",  -- ROS word 6a6
   "1000000000000000000000000000000101100000000100000000001100000000000000000000000000000000000100000000",  -- ROS word 6a7
   "0000001010000000000010000011011000000000000110010011010110000100000000000000000000000000110100110000",  -- ROS word 724
   "1000000000100000000111010000000101110000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 725
   "0000001010000000000010000011011000000000000110010011010110000100000000000000000000000000110100110000",  -- ROS word 726
   "0000001010000111100010000000000101110000000000010000011010000000011010000000000000010000010100000000",  -- ROS word 727
   "1000000000000000000000000000000101100000000100000000001100000000000000000000000000000000000100000000",  -- ROS word 7a4
   "1000000000000000000000000000000101100000000100000000001100000000000000000000000000000000000100000000",  -- ROS word 7a5
   "0000001010100000001101010000000000000000000000000100000000000011110010000000000000000100110100110000",  -- ROS word 7a6
   "1000001010000000000000000000000101100000000100000000001100000100000010000000000000000000110100110000",  -- ROS word 7a7
   "1000000000100000000111010000000101110000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 824
   "1000000000100000000111010000000101110000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 825
   "0000001010100000001101010000000000000000000000000100000000000011110010000000000000000100110100110000",  -- ROS word 826
   "1000001010000000000000000000000101100000000100000000001100000100000010000000000000000000110100110000",  -- ROS word 827
   "0000000000000010000000000000000000000000000000000000011100000000110000000000000000110000010000000000",  -- ROS word 8a4
   "0000000000000010000000000000000000000000000000000000011100000000110000000000000000110000010000000000",  -- ROS word 8a5
   "0000000000000010000000000000000000000000000000000000011100000000110000000000000000110000010000000000",  -- ROS word 8a6
   "0000000000000000000010000000000000000000000000000000011100000000110000000000000000000000000100000000",  -- ROS word 8a7
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 924
   "0000000000000000000000000010101000000000000000000011100001110000000000000000000000000100000100000000",  -- ROS word 925
   "1000000000000010100000000001000000000000000000000100101000000100010100000000000000000100000010110000",  -- ROS word 926
   "0000000000000000001010000010101000000000000000000011100000000000000000000000000000000000000100000000",  -- ROS word 927
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 9a4
   "0000000000000000000000000010101000000000000000010011010011110000000000000000000000000100000100000000",  -- ROS word 9a5
   "0000000000000010001010000000000000000001001000010011010010000100000010000000000000000000000100000000",  -- ROS word 9a6
   "1000000000000000000000000000000000000001011000010011010010000000000000000000000000000000000100000000",  -- ROS word 9a7
   "1000000000000010000000000000000000000000000000010100010100000010001001001000100000000100000001100000",  -- ROS word a24
   "0000000000000010000000000000000000000000000000010100010010000110001001001000100000000000000001100000",  -- ROS word a25
   "0000000000000010000000000000000000000000000000010100010100000110001001001000100000011000000000000000",  -- ROS word a26
   "0000000000000010000000000000000000000000000000010100010110000010001001001000100000011000000000000000",  -- ROS word a27
   "0000000000000000011100000000000000000000000000010101010010110100110111001111110000000110000100000000",  -- ROS word aa4
   "0011000000010000011101111000000000001000000000010101010100000000000010000000100001000100000100000000",  -- ROS word aa5
   "1000000000001000000000000000000000000000000000010101001010010100000000000000000000000000000100000000",  -- ROS word aa6
   "0011000000010000011101111000000000001000000000010101010100000000000010000000100001000100000100000000",  -- ROS word aa7
   "1000000000000000000000111000000000000000000010010110010010000101100000000000000000000000000100000000",  -- ROS word b24
   "1000001010000000000010000000000000000000000010110101001010000000000000000000000000000000000000001000",  -- ROS word b25
   "1000000000000111100000111000000000000000000101010110010010000001100000000000000000000000110100110000",  -- ROS word b26
   "1000001010000000000010000000000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word b27
   "0000000000000111000010000110100000000000000000010111010010000000000011101110100000000000000100000000",  -- ROS word ba4
   "0000001011000000000010000110100000000000000000010111000010000000000000000000001110000000000101000000",  -- ROS word ba5
   "0000000000000111100000000110111111010000000101010111010010000100000010000000000000000100110100110000",  -- ROS word ba6
   "1000000000000111000000000000000000000000000011010110100010000100000011001100000000000010000100000000",  -- ROS word ba7
   "1000000000010111100000000100101000000101010101011000001010000000000000000000000000000100110011100000",  -- ROS word c24
   "0000100000100000011000010101101000000010001000011000010000100000011001001111110000000111000111010000",  -- ROS word c25
   "0000000000000010000010000000000000001100001000011101011010000011111010000000000000000000000100000000",  -- ROS word c26
   "1000000000011111011100100001111000000101011000011001010010000000011000000000100001000000000100110000",  -- ROS word c27
   "0000000000010000000000000110011000010101010000011000011000001110100010000010110000000000000000000000",  -- ROS word ca4
   "0000000000000010000011000110101000001101001000011001010100000100000001001010100000000110000000110000",  -- ROS word ca5
   "1000000000000010000010110110111111100000000000011001010100000100000010000000000000000001011000000000",  -- ROS word ca6
   "1000000000000010000010110110111111100000000000011001010100000100000010000000000000000000001000000000",  -- ROS word ca7
   "0000110000100000000010000001111000000110100000011010010110000000000010000000000000000001000111010000",  -- ROS word d24
   "0000000000000010000000000001000000001100100000011011001010010100000000000000000000000100000101001000",  -- ROS word d25
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d26
   "1000110000100000000010000110010000000110110000011010010100000000000010000000000000000101000111010000",  -- ROS word d27
   "0000001010100000000010000000000000000101001100111011010000000100000000000000000000000100010001001000",  -- ROS word da4
   "0000000000001111000000000101111000000000000000011011010110000000000010000000000000000101011100001000",  -- ROS word da5
   "1000001011000000011100000111101000000000000000011010100000000100000010000011110000000100000001000000",  -- ROS word da6
   "0010100000000010000010000101111000001110010000011011001000000100000011010000100001000010000100001000",  -- ROS word da7
   "0000000000000011100000000001001000001100101001011100010100000100000010000000000000000100110100110000",  -- ROS word e24
   "0000001011001111010111000101101000000000000000111101010111010100000010000010100001110100000000000000",  -- ROS word e25
   "0000000000000000011110000100010010000000000000011100011100000000000010000000000000000000000100000000",  -- ROS word e26
   "1000001001101111000000000001000010000100010001011100011000000100000000000000000000000000000100000000",  -- ROS word e27
   "1000001010100000000010000111011001010101000000011001101000100000000010000000000000000000000001000000",  -- ROS word ea4
   "1000000000001111000010000101101001010000000000011001010110000100000010000000000000000100000100000000",  -- ROS word ea5
   "0000000000000010000000000000000000001100000000011100011110000100000010000000000000000000001000000000",  -- ROS word ea6
   "0000000001000000000000000000000001010000000000011111100000000110000100000000000000000000000011100000",  -- ROS word ea7
   "1000001010100000000010000000000000000110100000011111100100000001100100000000000000000101011101000000",  -- ROS word f24
   "0000000000000000000010000110101000000000000100111101101000000000000010000000000000000000000100000000",  -- ROS word f25
   "0000000000010010000010000000000000000100111000111110010100000010001000000000000000000000000100110000",  -- ROS word f26
   "0000000000000010010110010110011000001100000000111100011110000100000010000000100001000100000000001000",  -- ROS word f27
   "0000000000000010000000000000011000001110111000011111100110000110100010000000000000000100000100000000",  -- ROS word fa4
   "0001010000001010000010000000000000000000000000011111010010011000000000000000000000000000000100000000",  -- ROS word fa5
   "0000000000001001000010000000000000000000000000011111010110000100000000000000000000000000000100000000",  -- ROS word fa6
   "0000000011000111100000011001111000000000001000011111010100000000000000000000000000000000000011100000",  -- ROS word fa7
   "1000000000000010000010000001000000000011011000000011100000000100000010000000000000111000000000000000",  -- ROS word 028
   "1000000000000000000000000000000010000000000010001000100000000100000010000000000000000000000100000000",  -- ROS word 029
   "1000000000000000000000000001000000000000000000001111000010000000000000000000000000000000000100000000",  -- ROS word 02a
   "0000000000001111000010000000000000000000000000010000011100000000000010000000000000000000000100000000",  -- ROS word 02b
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a8
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0a9
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0aa
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0ab
   "0000000000000000000010000000000000000000000000001110000101111100000000000000000000000000000100000000",  -- ROS word 128
   "1000001011100000000000000000000000000001000000001110000001111100000000000000000000000100000011100000",  -- ROS word 129
   "1000001011100000000000000000000000000001000000001110000001111100000000000000000000000100000011100000",  -- ROS word 12a
   "1000001011100000000000000000000000000001000000001110000001111100000000000000000000000100000011100000",  -- ROS word 12b
   "1000000000100000000010000000000000000010000000000111100001111100000010000000000000000100000100000000",  -- ROS word 1a8
   "1000000000100111111100000000110000000001000000000111100011111100000010011101100000000000000101000000",  -- ROS word 1a9
   "1000000000100111111100000000110000000001000000000111100011111100000010011101100000000000000101000000",  -- ROS word 1aa
   "1000000000100111111100000000110000000001000000000111100011111100000010011101100000000000000101000000",  -- ROS word 1ab
   "0000000001001010000000000000000000000000000101100100010110000100000010000000000000000000000001000101",  -- ROS word 228
   "1000000001000000000010000110001000000000000000000111011010000000000000000000000000000100000100000011",  -- ROS word 229
   "1000000001001010000000000000000000000000000101100100010110000100000010000000000000000000000100000101",  -- ROS word 22a
   "0000000000000000000011100000000011110000000000000111010010000100101000000000000100000100010011010000",  -- ROS word 22b
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a8
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2a9
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2aa
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2ab
   "1000000000000100100010000000000000000000000110100110001000000000000000000000000000000100000100000000",  -- ROS word 328
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 329
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 32a
   "0000000000000100100010000000000000000000000110100100101000000000000010000000000000000000000100000000",  -- ROS word 32b
   "0000000000000000000010000000000000000000000000000111010110000000000010000000000000000000000100000000",  -- ROS word 3a8
   "1000000000000000000010000000000000000000000000000111010110000000010010000000000000000100000100000000",  -- ROS word 3a9
   "1000000000000000000010000000000000000000000000000111010110000100110100000000000000000100000100000000",  -- ROS word 3aa
   "1000000000000000000010000000000000000000000000000111010110000000010010000000000000000100000100000000",  -- ROS word 3ab
   "0000000000000011000000000101000000000001011000010010010010000000111001001100000000000011000000000000",  -- ROS word 428
   "0000000000000000000011000111011000000000000000001110010110000111110110000000000000000000000100000000",  -- ROS word 429
   "0000000100000010011110000001011000000001001000001000010100000011011111001110111010000011110100000000",  -- ROS word 42a
   "1000000000000011000000000101000000000001011000010010010010000000000000000000100000000100000000110000",  -- ROS word 42b
   "0000001000000000000000000110000000000011011000001001010100000000001111110000101010000000000011100000",  -- ROS word 4a8
   "0000000000010010000000000000000000000011010000001100001010010100000100000000001010000001001001000000",  -- ROS word 4a9
   "0000000000000000000000000111000000000000000000001001010100000000000000000000000000000100000100000000",  -- ROS word 4aa
   "0000000000000111100010000000000000000000000000110001100110000001000010000000000000000100100000110000",  -- ROS word 4ab
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 528
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 529
   "0000001001000000000010000000000000000000000001010011000000000000000010000000000000000000000100000000",  -- ROS word 52a
   "1000000000000000000010000000000000000000000000010000001110000001100000000000000000000100000100000000",  -- ROS word 52b
   "0000000000000111000000110110000000000000000011010010001101001100001111111011000000000100000100000000",  -- ROS word 5a8
   "1000000000000111000000110110000000000000000011010010001101001100001111111001000000000100000000000000",  -- ROS word 5a9
   "0000000000001010000001100000000110010000000101100000010100000000000010000000000000000100000100000000",  -- ROS word 5aa
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 5ab
   "1000000000000000000010000000000000000000000000001100011000010100000000000000000000000100000100000000",  -- ROS word 628
   "0000000000100000000010000111111000000011010000010001011000000000000010000000000000000000000100000000",  -- ROS word 629
   "0000000000000000000010000101101000000000000000001111001110000000000000000000000000000000000100000000",  -- ROS word 62a
   "1000000000000000000010011000000000000000000101101101010100000000000000000000000000110100000100000011",  -- ROS word 62b
   "0000000000000000000010000000000000000000000010001101010100000000000010000000000000000000000100000000",  -- ROS word 6a8
   "1000000000100000000010000000000000000011010000010001011000000001100000000000000000000100000100000000",  -- ROS word 6a9
   "1000000000000111100010000000000000000000000000101010010110000100110100000000000000000100110100110000",  -- ROS word 6aa
   "1000001001001001100000000000001011010000000000110000010100000100000000000000000000000000000100000000",  -- ROS word 6ab
   "0000001001000000000010000000000000000000000000101110000110000101010010000000000000000100000000000010",  -- ROS word 728
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 729
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 72a
   "1000000000001001000000000101001000000000000000001101010100000100000010000000000000000000000100000000",  -- ROS word 72b
   "1000000000000000000010000000000000000000000101001111010100000100000010000000000000000100000100000000",  -- ROS word 7a8
   "1000000000000000000011011101010000000000000000010000010101010100000010000000000000000000000011100000",  -- ROS word 7a9
   "0000000000010010000000000000000000000011010000101011010100000100000000000000000000000001011000000000",  -- ROS word 7aa
   "0000000000001010000000000011010000000000000001001111010100000000000010000000000000000100000100000000",  -- ROS word 7ab
   "1000000000000111100010000101110000000000000000001100010010001100011110000000000000000100110100110000",  -- ROS word 828
   "0000000000000000000001010000000010000000000000010001011110000000000000000000000000000100000100000000",  -- ROS word 829
   "0000001010000011100010000000000101100000000101001011001010000000000010000000000000000101011000000000",  -- ROS word 82a
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 82b
   "1000000000001010100000000000000000000001111000010000010010111000011110000000000000000101011000000000",  -- ROS word 8a8
   "0000000001100000000010000000000000000010010000000000011110000000000010000000000000000001011111100000",  -- ROS word 8a9
   "0000000000001010100000000000000000000001111000001111010010111000011110000000000000000001011000000000",  -- ROS word 8aa
   "0000000000010111100010000101100110010011010101001110010100000100000010000000000000000000000100000000",  -- ROS word 8ab
   "0000000000000000010110000000000000000000000000000111010010000001101010000000000000000000000100000000",  -- ROS word 928
   "1000000000000010010110000000000001000000000001000011101000000100000010000000000010000000000000000000",  -- ROS word 929
   "0000001011000000000000111110100000000000000011001111010001001000000000000000000000000000000001000000",  -- ROS word 92a
   "0000000001000000000000111110100000000000000011001111010001001000000000000000000000000000000011100000",  -- ROS word 92b
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9a8
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9a9
   "1000000000000000000010000000000000000000000000010000001110000000000000000000000000000100000100000000",  -- ROS word 9aa
   "0000000000000000000010000000000000000000000000010010011000000000000010000000000000000000000100000000",  -- ROS word 9ab
   "1000000000000000000000000010000000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word a28
   "0000000000000010000000000000000000000000000000010100010100000110001001001000100000011000000000000000",  -- ROS word a29
   "1000000000000000000000000010000000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word a2a
   "0000000000000010000000000000000000000000000000010100010110000110001000000000000000000100000101100000",  -- ROS word a2b
   "1000000000000000011110010000000000000000000000010101101010000000000000000011100001000100000100000000",  -- ROS word aa8
   "0000000000000000011100000000000000000000000001010101010101000100110111001111110000000110000100000000",  -- ROS word aa9
   "1000000000000000011110010000000000000000000000010101101010000000000000000011100001000100000100000000",  -- ROS word aaa
   "1000000000001000000000000000000000000000000000010101001010010100000000000000000000000000000100000000",  -- ROS word aab
   "0000000000000000011110000111101000000000000000010110010100000101010111001110110000000110000000000000",  -- ROS word b28
   "1000000000000000000010000000000000000000000000010110001000000100000011010000100000000110000100000000",  -- ROS word b29
   "1000001001001110111100000000000000000000000000010110010100000000000011001110110000000110000000000000",  -- ROS word b2a
   "1000001001000101000000000101001000000000000000010110001110000000000010000000000000000000000100000000",  -- ROS word b2b
   "1000000000000111000010000110111000000000000000010111001010000100000001001100000000000000000000000000",  -- ROS word ba8
   "1000000000000111000000000110000000000000000000010111010100000100000000000000000000000000000100000000",  -- ROS word ba9
   "1000000000000111000010000110010000000000000000010111010100000100000011101110100000000100000100000000",  -- ROS word baa
   "1000000000000000011110000111011000000000000000010111010110000000000000111100000000000010000000000000",  -- ROS word bab
   "0000000000000010000000000000000000000001111000011111010000000000000000000000000000000100000100110000",  -- ROS word c28
   "0000000000010010000000000000000000000110010000011001011100000100000000000000000000000001000000000000",  -- ROS word c29
   "1000001001000000011100000001111000000000000000011000000100000100010101110100000000000110000000000000",  -- ROS word c2a
   "1000000001110000011110000110011000000101000000011001000000000000010101110100000000000010110000110000",  -- ROS word c2b
   "1000000001000010010110000110110000000000000000011001010110000100000000000000000000000000001000000000",  -- ROS word ca8
   "0000000001000010010110000110110000000000000000011001010110000100000000000000000100000000001100000000",  -- ROS word ca9
   "0000001101000000011110110110101000000000000000011001010010000110001000000000100000000100000000000000",  -- ROS word caa
   "0000000110000000000010110110110111100000000000011001010110000000000001001010000100000110000000000000",  -- ROS word cab
   "1000001010010000011111000101101000000101010000011010001110000100000000000000100001000000000001000000",  -- ROS word d28
   "0000100000100000000000000000000000000110111000011010010100000100011000000000000000000101000111010000",  -- ROS word d29
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d2a
   "1000110000000000000010000000000000000000000000011011001010100000000010000000000000000101000111010000",  -- ROS word d2b
   "0010100001000000000000000110101000000000000000011011010100000100000001010000100001000010000000110000",  -- ROS word da8
   "1000000000000010000010000000000000001100111011011011100100000100000000000000000000000000010001001000",  -- ROS word da9
   "0000000000000010011100100110101000000000000000011011010110000110001000000000100001000101101101000000",  -- ROS word daa
   "1000000001000111000010000000000000000000000000011011011000000110001000000000000000000001101000110000",  -- ROS word dab
   "1000001010000000000000000010111011010000000100011101011000000100000010000000000000010000010100000000",  -- ROS word e28
   "1000001010000000000010000010111000001100110100111100010010000010001010000000000000010100010100101000",  -- ROS word e29
   "0000001010000010000000000000000000000000000000011100000000000000000010000000000000000101000111100000",  -- ROS word e2a
   "1001010000000000000010110000000000000000000111011100010110000100000000000000000000000100000100000000",  -- ROS word e2b
   "0000001010000010000000010000000000001100100000011100101010000011111010000000000000010100010100000000",  -- ROS word ea8
   "1000000000000010000000000000000000001100000000111100011110000100000010000000000000000100000000001000",  -- ROS word ea9
   "0000001010000010000010000000000000001100100000011100011110000011111010000000000000010000010100000000",  -- ROS word eaa
   "1000000000000010000000000101101000001100011000011101010110000000000000000000000000000000000100110000",  -- ROS word eab
   "1000000001000000010110001000000000000000000000011110010110000000000001010000100001000010000000000000",  -- ROS word f28
   "0000000000000111100010000101110000001100011101011110010100000100011010000000000000000100000001000000",  -- ROS word f29
   "1000001010000000000010000110101000000000000000111101101000000000000000000000000000000000010001001000",  -- ROS word f2a
   "1000001010000000000010000010111000000000000000011110010010000000000010000000000000000000010001001000",  -- ROS word f2b
   "1000001010001111000010000000000000000000000000011111011000000000000000000000000000000000000001000000",  -- ROS word fa8
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fa9
   "1000001010000011100000000000000000000011011000011111011110000000000010000000000000111100000000000000",  -- ROS word faa
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fab
   "1000000000100000000000000000000000000101000000000000001010000000000010000000000000000000000100000000",  -- ROS word 02c
   "0000001010000000000000000010000000000000000000000000001000000000000000000000000000000000000001000000",  -- ROS word 02d
   "0000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 02e
   "1000001010000000000000000000000101100000000101000001101000000100000010000000000000000000110100110000",  -- ROS word 02f
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0ac
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0ad
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0ae
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0af
   "0000001011010000000001000111011000000001000000001110000001111100000010000000000000000000000011100000",  -- ROS word 12c
   "0000001011100000000000000000000000000001000000001110000111111100000010000000000000000000000011100000",  -- ROS word 12d
   "1000001011100000000000000000000000000001000000001110000001111100000000000000000000000100000011100000",  -- ROS word 12e
   "1000001011100000000000000000000000000001000000001110000001111100000000000000000000000100000011100000",  -- ROS word 12f
   "0000000000100111111100000000110000000010000000000011100101111100000011111101100000000100000111100000",  -- ROS word 1ac
   "1000000000100111111100000000110000000001000000000001100011111100000010011101100000000000000111100000",  -- ROS word 1ad
   "1000000000100111111100000000110000000001000000000111100011111100000010011101100000000000000101000000",  -- ROS word 1ae
   "1000000000100111111100000000110000000001000000000111100011111100000010011101100000000000000101000000",  -- ROS word 1af
   "0000000001001010000000000000000000000000000101100100010100000100000010000000000000000100000101000100",  -- ROS word 22c
   "1000000000000000000010000000000000000000000000000111011010000000010010000000000000000100010100100000",  -- ROS word 22d
   "1000000001001010000000000000000000000000000101100100010100000100000010000000000000000100000000000100",  -- ROS word 22e
   "0000000000000000000010000000000011110000000000000111010010000100101000000000000100000100010011010000",  -- ROS word 22f
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2ac
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2ad
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2ae
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2af
   "0000000000000000001000000000000000000000000000000110010100000100000010000000000000000100000100000000",  -- ROS word 32c
   "0001010000000000000010000000000000000000000110100100101000000000000010000000000000000000000100000000",  -- ROS word 32d
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 32e
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 32f
   "0000001001000000000010000000000110000000000000000110000000000011001110000000000000000000000100000000",  -- ROS word 3ac
   "0000001001000000000010000000000110000000000000001000000000000011001100000000000000000000000100000000",  -- ROS word 3ad
   "1000001001000000000010000000000110000000000000001000000000000100000000000000000000000100000100000000",  -- ROS word 3ae
   "1000001001000100100010000000000110000000000000001100010100000100000010000000000000000100000100000000",  -- ROS word 3af
   "0000000000000000001000000000000000000000000000101011001000000000000010000000000000000100000100000000",  -- ROS word 42c
   "1000000000000000000000000000000011010000000000010101001010000000000000000000000000000000000100000000",  -- ROS word 42d
   "0000001011000000000000111110100000000000000011010001010001001000000000000000000000000000000001000000",  -- ROS word 42e
   "0000000001000000000000111110100000000000000011010001010001001000000000000000000000000000000011100000",  -- ROS word 42f
   "1000000000000110000000110110001000000000000000001111101001001100001111101100000000000100000000100000",  -- ROS word 4ac
   "1000000000000110000000101110010000000000000011001111001000001100000010000000000000000100000000100000",  -- ROS word 4ad
   "1000001011000000000000111110100000000000000011010011010001001000000000000000000000000100000001000000",  -- ROS word 4ae
   "1000000001000000000000111110100000000000000011010011010001001000000000000000000000000100000011100000",  -- ROS word 4af
   "1000001011000000000010100110000000000000000011001010000000000011000100000000000000000000000001000000",  -- ROS word 52c
   "1000000001000000000010100110000000000000000011001010000000000011000100000000000000000000000011100000",  -- ROS word 52d
   "1000001001000100100010000000000000000000000000001010010010000000000000000000000000000100000100000000",  -- ROS word 52e
   "1000001001000100100010011000000000000000000101101101010100000000000000000000000000110100000100000011",  -- ROS word 52f
   "0000000000100000000000000111000001010011010000001011010110000000000010000000001000000000000000000000",  -- ROS word 5ac
   "1000000000000111000000000000000000000011011000001000100010000100000011100000101000000000000100000000",  -- ROS word 5ad
   "1000001011000000000000111110100000000000000011001001010011001000000000000000000000000100000001000000",  -- ROS word 5ae
   "1000000001000000000000111110100000000000000011001001010011001000000000000000000000000100000011100000",  -- ROS word 5af
   "0000000000010010000000000111000011010011010000001101101010000000000010000000001010000000000001000000",  -- ROS word 62c
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 62d
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 62e
   "1000000000000000000010000000000001100000000000010001001100000100000010000000000000000100000100000000",  -- ROS word 62f
   "1000000000000111000000000000000000000011011000001101010110000000000011100000101000000000000100000000",  -- ROS word 6ac
   "1000000000010010000000000110011000000011010000001110010110000000000000000000001000000100000000000000",  -- ROS word 6ad
   "0000000101000000011100110000000111100000000000000010100100000000000011001110000100000110101100000000",  -- ROS word 6ae
   "1000000000000000000001000000000000000000000000000011100010000000000010000000000000000000000100000000",  -- ROS word 6af
   "1000000000000000011010000000000000000000000000001001000010000100000010000011100000000000000000000000",  -- ROS word 72c
   "1000000000100000000000000111000001010011010000001101010110000000000000000000001000000100000000000000",  -- ROS word 72d
   "1000001001000010000000000110011000000000000000001010011000011000000010000000000000000000000100000000",  -- ROS word 72e
   "0000000000001101000000000000000000000000000000000011011110000000000000000000000000000100000100000000",  -- ROS word 72f
   "0000000000000111000000000000000000000000000011001000100010000100000011001100001000000010000000000000",  -- ROS word 7ac
   "1000000000000111000000000000000000000000000011001011010110000000000001001100001000000110000000000000",  -- ROS word 7ad
   "1000001001000000000010000000000000000000000000001100011110000000000000000000000000000100000100000000",  -- ROS word 7ae
   "0000000001000100100000000110011000000000000000001101011110000000000000000000000000000000000001000000",  -- ROS word 7af
   "1000000000000111000000000000000000000000000000010010101000000100000001001100000000000010000100000000",  -- ROS word 82c
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 82d
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 82e
   "0000000000000000000010000000000001100000000000100000001110000000000010000000000000000000000100000000",  -- ROS word 82f
   "1000000000000000000010000000000000000000000000010111000100000100110110000000000000000100000100000000",  -- ROS word 8ac
   "1000000000000000000010000000000000000000000000000110011110000101000110000000000000000100000100000000",  -- ROS word 8ad
   "0000000000100000001101010000000000000000000000000100000000000011110010000000000000000100000100000000",  -- ROS word 8ae
   "0000001010000000000010000011011000000000000000010010010110000100000010000000000000010000010100000000",  -- ROS word 8af
   "0000000000000000000010000000000000000000000000010011101000000000000011101000000000000100000000000000",  -- ROS word 92c
   "0000000000100000000010000000000000000011010000001001001100000100010100000000000000000000000100000000",  -- ROS word 92d
   "0000000000000011000000000101000000000001011000000100101000000111011111001100000000000110000100110000",  -- ROS word 92e
   "0000000000001010000010000000000000000000000000010011101010000100000000000000000000000000000100000000",  -- ROS word 92f
   "1000001001000000000000000001110000000000000000010010010110000000000000000000000000000000000100000000",  -- ROS word 9ac
   "1000001001000000000000000001110000000000000000010010010110000000011100000000000000000100000011100000",  -- ROS word 9ad
   "0000000000001010000000000100110010010000000000010001010110000100011110000000000000000100000100000000",  -- ROS word 9ae
   "0000000001001010000010000100110010010000000000010010011110000000000000000000000000000100000011100000",  -- ROS word 9af
   "0000000000000010000000000000000000000000000000010100010110000110001000000000000000000100000101100000",  -- ROS word a2c
   "1000000000000010000000000000000000000000000000010100010110000100000010000000000000000000000101100000",  -- ROS word a2d
   "1000000000000000000000000010000000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word a2e
   "0000000001100000000010000110010000000001110000010100011000000000000000000000000000011100110011100000",  -- ROS word a2f
   "0000000000000000000010000011010000000000010000010101001010000000000000000000000000000000000100000000",  -- ROS word aac
   "1000000000000111100010000000000000000000000101110101100110000100000010000000000000000000000011100000",  -- ROS word aad
   "0000000000000000000010000101101000000000000000010101010111111100000000000000000000000000000100000000",  -- ROS word aae
   "0000000000000000000010000101101000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word aaf
   "1000000000000000000010000100000011010000000000000000000001100000000000000000000000000100000100000000",  -- ROS word b2c
   "1000000000000111100000000101001000000000000001110110001110000100000000000000000000000000110100110000",  -- ROS word b2d
   "1000000000010010000010000000000000010011010000110110010110000100000010000000000010000000000000000000",  -- ROS word b2e
   "0000000000000000000010000000000000000000000101010110011000000000000000000000000000000000000100000000",  -- ROS word b2f
   "1000000000000111000000000000000000000000000000010111010110000000000011000100110000000110000000000000",  -- ROS word bac
   "0000000000000010000000000000000000000000000000010111010110000100000000000000001110000100000111100000",  -- ROS word bad
   "0000000000000010011110000000000000000000000000010111010110000100000010000000100000000000000101000000",  -- ROS word bae
   "0000000000000111000000000000000000000000000000010111011100000100000001001100000000000110000100000000",  -- ROS word baf
   "0000000000001111011100000000000000000000000000011000001010111100000010000000100000000000110000110000",  -- ROS word c2c
   "0000000000000010000000000110011000000000000000011000010010000000000000000000000000000100110100110000",  -- ROS word c2d
   "0000001010000000000010000000000000000000000000011001100100000100011010000000000000000000010111010000",  -- ROS word c2e
   "1000000000000010000000000000000000001100110000011001101000000000000000000000000000000001011111100000",  -- ROS word c2f
   "0000000110000000011010011110110111100000000000011001010100000010001000000011100101000000001100000000",  -- ROS word cac
   "1000000000000000000001000110101000000000000000011001010100000100000001001010100000000110000000000000",  -- ROS word cad
   "0000000011000111011110000110011000000000000000011001011110010100000001001000100000000010000110001000",  -- ROS word cae
   "0000000000000010010110000000000000000010011000011100011000000000000011000110110000000110010000000000",  -- ROS word caf
   "0000000001000000000000110000000001010000000111011010011110000000000000000000000000000100110100110000",  -- ROS word d2c
   "0000100000100000000000000111011000000110101000011010010010000100011000000000000000000101000111010000",  -- ROS word d2d
   "1000000000000000011111000110110000000000000000011011000000000000000000000000100001000100000100000000",  -- ROS word d2e
   "0000000000000000011101100110110000000000000000011011000000000000000000000000100001000100000100000000",  -- ROS word d2f
   "1000000000100111100010000110110000000101001101011011010000000000000010000000000000000100010111100000",  -- ROS word dac
   "0011100001000111000000000001111000000000000000011011011000000100000010000000100101000100001100000000",  -- ROS word dad
   "1010101011000000000000000000000000000000000000011011010100000100000011010000100001000110000000000000",  -- ROS word dae
   "1000000000000000000010000101011000000000000000011011010110000000000000000000000000011001101001001000",  -- ROS word daf
   "0000000000000010000010000000000000001100100000011100010110000000000010000000000000000001000111010000",  -- ROS word e2c
   "1000000000100000000010000000000000000100000000011111001010000100000000000000000000000100000100000000",  -- ROS word e2d
   "0000000000000000000010000000000000000000000010011100010110000100000010000000000000000000000100101000",  -- ROS word e2e
   "1000000001000000000010010000000000000000000000011100011000000000000000000000000000110001011000000000",  -- ROS word e2f
   "1000000000011111000010000110011000000011010000011101010010000000000000000000000000000100000100000000",  -- ROS word eac
   "0001010000000111100010110000000000000000000000111101010110000100000000000000000000000000110100110000",  -- ROS word ead
   "1000000000000000000010000001001000000000000000011101001110000000000010000000000000000100000100101000",  -- ROS word eae
   "1000000000000010000000000000000001011100110000011101001110000100000000000000000000000100000001000000",  -- ROS word eaf
   "1000000000000000011010000110011000000000000000011110011100000100000000000000000000000100000100000000",  -- ROS word f2c
   "0000000000001111000000000000000000001100010000011110010110000100000000000000000000000100000100000000",  -- ROS word f2d
   "1000000000000010000010000000000000001100001100111110010110000100000010000000000000000000001000000000",  -- ROS word f2e
   "1000000001000000000010000000000000001110110000011110100110000100000000000000000000000100000100110000",  -- ROS word f2f
   "0000000000000000000010110000000111100000000000011111010111001100000000000000000000000000000100000000",  -- ROS word fac
   "0000000000000000000010000000000000000000000001011111010010000000000010000000000000000000000100000000",  -- ROS word fad
   "0011110000000000000010000000000000000000011000011111010010000100000010000000000000000000000100000000",  -- ROS word fae
   "0000000000011011100010000000000000001011101000011111011010000100000000000000001110000000000100001000",  -- ROS word faf
   "0000000000000000000010000000000011110000000000000011000000000011001110000000000000000000000100000000",  -- ROS word 030
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 031
   "0000000000000000000000000000001011110000000101000010000000000011001110000000000000000100000100000000",  -- ROS word 032
   "1000000000000111000000000000000001100000000000101000001110000000000000000000000000000000000100000000",  -- ROS word 033
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b0
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b1
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b2
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b3
   "1000000000000000000000000011010000000000000011110011010011111100000000000000000100000000010110100000",  -- ROS word 130
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 131
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 132
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 133
   "0000000000000111101010000000010000000000000000000100100001111100000010000000000000000100000011100000",  -- ROS word 1b0
   "0000000000000111101010000000010000000000000000000100100001111100000010000000000000000100000011100000",  -- ROS word 1b1
   "0000000000000111101010000000010000000000000000000100100001111100000010000000000000000100000011100000",  -- ROS word 1b2
   "0000000000000111101010000000010000000000000000000100100001111100000010000000000000000100000011100000",  -- ROS word 1b3
   "0000000000000111100010000100110100110000000000000100000101100100000010000000000000000100000011100110",  -- ROS word 230
   "1000000000000111100010000100110100000000000000000100000111100100000010000000000000000000000011100101",  -- ROS word 231
   "0000000000000111100000000000001100010000000000000111000111100100000000000000000000000100000111100100",  -- ROS word 232
   "1000000000000111100000000000001100100000000000000111000111100100000010000000000000000000000111100111",  -- ROS word 233
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2b0
   "0000001010000100111110000101111000000000000100000111001100000100000000000000000000000000000111100001",  -- ROS word 2b1
   "0000001010000100111110000101111000000000000100000111001100000100000000000000000000000000000111100001",  -- ROS word 2b2
   "1000001010000100111110000101111000000000000100000111001100000000000000000000000000000100000111100001",  -- ROS word 2b3
   "1000001001000000011100000000000000000000000001000111000010000000000000000000000000000000000100000000",  -- ROS word 330
   "1000000000000111000010101110010000000000000011001000101000001100000010111100110000000100000100000000",  -- ROS word 331
   "0000000000000111000000000000000000000000000000001010010110000010001110110100000000000000000000000000",  -- ROS word 332
   "0000000000000111000000000000000000000000000000001011100110000110001110110100000000000000000000000000",  -- ROS word 333
   "0000001010000010000010000000001000000000000000000101000000000011001110000000000000000000000101000111",  -- ROS word 3b0
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 3b1
   "1000001010000010000010000000001000000000000000000101000000000011001110000000000000000000000000000111",  -- ROS word 3b2
   "1000000000000111000010000001001101100000000000100000001110000000000000000000000000000100000100000000",  -- ROS word 3b3
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 430
   "0000000000000111000010101110010000000000000011001000101000001100000000111100110000000000000100000000",  -- ROS word 431
   "0000000000000111000010100110000000000000000011001010000100000011000100110100000000000100000000000000",  -- ROS word 432
   "1000000000000111000010100110000000000000000011001001100100000011000100110100000000000000000000000000",  -- ROS word 433
   "1000000000000111000010101110010000000000000011001001011000001100000001110000100000000100000100000000",  -- ROS word 4b0
   "0000000000000000000010000000000000000000000000001101001110100000000000000000000000000000000100000000",  -- ROS word 4b1
   "1000000000000000000010000000000000000000000101101001001110010000000100000000000000000100000100000000",  -- ROS word 4b2
   "1000000000000000000000000001001101100000000000100000001110000000000010000000000000000000000100000000",  -- ROS word 4b3
   "0000000000000111000010101110010000000000000011001010011000001100000001100000100000000100000000000000",  -- ROS word 530
   "1000000000000111100010110000000111100000000000001010011100000000000000000000000000000001000000000000",  -- ROS word 531
   "1000000000000000000000000000000101100000000101100000010010010000000010000000000000000000000100000000",  -- ROS word 532
   "0000001011000111100000110000000111100000000000001010011100000000000000000000000000000001011000000000",  -- ROS word 533
   "1000000000000010000000000000000000000011011000001011011000000000000010000000000000111100000000000000",  -- ROS word 5b0
   "1000000000010111100010000000000000000011010101001011011010000100000010000000000000000100110100110000",  -- ROS word 5b1
   "0000000000000000000010000000000000000000000000001111011000000100000000000000000000000000000100000000",  -- ROS word 5b2
   "0000000000000000000010000000000000000000000000000101101000000011111000000000000000000000000100000000",  -- ROS word 5b3
   "0000000000000100100010000000000110000000000000001000000000000011001100000000000000000000000100000000",  -- ROS word 630
   "1000000000000111000010000011010000000000000000001111010100000010001001011000100000000100000100000000",  -- ROS word 631
   "0000000000000100100000000001000110000000000000001111000100000000000010000000000000000100000100000000",  -- ROS word 632
   "0000000000000111000010000011010000000000000000001111010100000010001001001100000000000100000000000000",  -- ROS word 633
   "0000000000000000000000000101001000000000000000010001100010000000000000000000000000000100000100000000",  -- ROS word 6b0
   "0000000000000000000010000000000000000000000000000000010110000100000010000000000000000000000100000000",  -- ROS word 6b1
   "0000000000000000000010000000000000000000000000010000100000000011011100000000000000000000000100000000",  -- ROS word 6b2
   "0000000000000000010000000000000000000000000000010000001110000100000010000000000000000100000100000000",  -- ROS word 6b3
   "1000000000000000000010011101111000000001101000000001101010000000000010000000000000000001000000000000",  -- ROS word 730
   "0000000000000000000010011101111001010001101000000001101010000000000000000000000000000101000000000000",  -- ROS word 731
   "0000000000000000000010000000000000000000000010001000010110000000000000000000000000000000000100000000",  -- ROS word 732
   "0000000000000000011000000000111000000000000000000100101000000000000000000000000010000000000000000000",  -- ROS word 733
   "1000000000000000000000000001000000000000000101001011011100000100000000000000000000000000000100000000",  -- ROS word 7b0
   "0000000000000000000010000000000000000000000101001011011100000100000000000000000000000000000100000000",  -- ROS word 7b1
   "0000000000000010000000000000000000000000000000000000001001100000000000000000000000111000000000000000",  -- ROS word 7b2
   "1000000000000000000010000000000000000000000001001110011000000100000010000000000000000100000100000000",  -- ROS word 7b3
   "0000000000000000000010000111100000000000000000001011000010000100000000000000000000000000000100000000",  -- ROS word 830
   "0000001010000000000010000110010101100000000100001111000100000100000000000000000000010000010100000000",  -- ROS word 831
   "0000000000000000000010000000000000000000000000010000011100000110001000000000000000000000000100000000",  -- ROS word 832
   "0000000000001110100010000000000000000000000001001111011000000100000010000000000000000000000100000000",  -- ROS word 833
   "0000001010000000000010000000000000000000000100001101010100000100000000000000000000010000010100000000",  -- ROS word 8b0
   "1000001010000000000010000101101101110000000000000000001000000000000000000000000000000000000011100000",  -- ROS word 8b1
   "0000000000001001011110011101111000000000000000010001000100000100001010000010110000000100000000110000",  -- ROS word 8b2
   "0000000000000000000010000000101000000000000000010000011000000100000010000000000000000000000100000000",  -- ROS word 8b3
   "1000000000000111100010000000000000000000000000001010010010000000000000000000000000000100110100110000",  -- ROS word 930
   "0000000000100000000010000000000000000011010000010001011000000000000010000000000000000000000100000000",  -- ROS word 931
   "0000000000000000000010000110110000000000000000010010011100000100000010000000000000000000000100000000",  -- ROS word 932
   "1000000000000111100010000000000000000000000101010010011010000100000000000000000000000100110100110000",  -- ROS word 933
   "0000000000000000000010000000000000000000000110110011011000000000000010000000000000000000000100000000",  -- ROS word 9b0
   "1000000000000000000010000000000000000000000000101110000000000100000010000000000000000100000100000000",  -- ROS word 9b1
   "1000000000001110001010000000000000000000000000001000100000000100000010000000000000000100000100000000",  -- ROS word 9b2
   "0000001010000001100000000000000101100000000100001011001010000000000010000000000000000000000011100000",  -- ROS word 9b3
   "1000000001000111111110000110110000000000000000010100011000000000000010000000110000011001011000000000",  -- ROS word a30
   "1000000001000110000000000000000000000000000000010100011000000100000000111100110000011011011100110000",  -- ROS word a31
   "0000000000000000000000000000000010000000000000110100011010000000000000000000000000011100000100000000",  -- ROS word a32
   "1000000000000000000010000101101000000000000000010100011100000000000000000000000000000000000011100000",  -- ROS word a33
   "0000001010000000000000000010000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word ab0
   "1000000000000000000010000000000000000000000101010110000011000000000010000000000000000100000100000000",  -- ROS word ab1
   "0000000000000000000010000000101000000000000101010101011101000000000000000000000000000000000100110000",  -- ROS word ab2
   "1000000000000000000010000000000000000000000000010101011010000000101110000000000000000100000100000000",  -- ROS word ab3
   "0000000000000000000000000000000011010000000010011111101000000000101110000000000000000100000100000000",  -- ROS word b30
   "0000000000010111100000000000000000000010111000010111100000000000000010000000000000000100110100110000",  -- ROS word b31
   "0000000000000010000000000000000000000011011010010110011010000100000010000000000000000000000000001000",  -- ROS word b32
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word b33
   "1000000000000000010010000011010000000000000000010111011010000100000000000000000100000100010110100000",  -- ROS word bb0
   "0000000000000000000000000011010000000000000001010111011010000000000000000000000100000100010110100000",  -- ROS word bb1
   "0000000000000000010000000000000000000000000000010111011010000100000000000000000000000100000100000000",  -- ROS word bb2
   "0000000000000000000000000001101000000000000000001000100000000100000010000000000000000100000100000000",  -- ROS word bb3
   "0000000000000010000011000001111000001101010000011000011010000100000010000000000000111001011100000000",  -- ROS word c30
   "0000000000000111100000000100101000000000000101011000001010000000000000000000000000000100110100110000",  -- ROS word c31
   "0000000000000111100000000100101000000000000101011000001010000000000000000000000000000100110100110000",  -- ROS word c32
   "1000000001010000000000000000011000000101100000011000011000000000000000000000000000000100000001000000",  -- ROS word c33
   "0000000000010010000001000101101000000101101000011001001000000011001000000000000000000001011000000000",  -- ROS word cb0
   "1000000000010010000011000000000010000101101000011001001000000100000000000000000000000001011000000000",  -- ROS word cb1
   "0000001101000000011110011000000000000000000000011001011000000100000010110100001110000010100100000000",  -- ROS word cb2
   "1000000000010111000010011110110000000101000000011001011010000000000001001100000000000100000100001011",  -- ROS word cb3
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d30
   "1000000001010000011110100001001000000101011000011001010110000000000010000000100001000000000001000000",  -- ROS word d31
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d32
   "1000000000010010000000000001000000000100001000011010011010000000000000000000000000000101000000000000",  -- ROS word d33
   "0000000000000110000011100110010000001101011000011011011010000000000000000010100001000000000111100000",  -- ROS word db0
   "1000000000000111000000000000000000000000000101011010011100000000000001001100000000000100000000000000",  -- ROS word db1
   "0000000000000010011100000100011010001100111000011101010110000000000000000000000000000000010000000000",  -- ROS word db2
   "1000000000000000000000000111101000000000000011011011011000000000000010000000000000000000000100000000",  -- ROS word db3
   "0000000000010010000000000000000000000100110000011100010100000011111010000000000000000000010000000000",  -- ROS word e30
   "1000000000100000000000011000000000000110011000011001011010000100000000000000000000000000000100000000",  -- ROS word e31
   "0000001010000000000010000010111000000000000100111100011000000100000010000000000000000001101111100000",  -- ROS word e32
   "0000000000000010000010111100000000001100111000111101001100000000000011010000100001000101101000110000",  -- ROS word e33
   "0000000000001011100010000000000000000000000000011101100110000100000010000000000000000000000100000000",  -- ROS word eb0
   "1000000000000111111010000000000000000000000101011101011000000100000000111100000000000010110000110000",  -- ROS word eb1
   "0000000000101011100000000000000000000101011011111101011100000010001000000000000000000100000100000000",  -- ROS word eb2
   "0000000000000010000000011000011000000000000000011100001010000000000010000000000000000100000100101000",  -- ROS word eb3
   "0000000000001111000010000000000000000000000000011110100010000000000000000000000000000100000000001011",  -- ROS word f30
   "1000000000001111000010000000000000000000000100111110011000000100000000000000000000000000000000001011",  -- ROS word f31
   "0000000000000000000010000000000000000000000001011110100100000000000000000000000000000000000100000000",  -- ROS word f32
   "0000000001000000000010000000000000001100100000011111001000000011111011101100000000000111011000001000",  -- ROS word f33
   "1000000000001011000010100110101000000011101000011111011000000001001111001100000000000001000001110000",  -- ROS word fb0
   "1000001101000000000010000110011000001110110000011111011000000100000000000000000100000101011100000000",  -- ROS word fb1
   "1000000000000000011110100110110000000000000000011111011000000100101110000000100000000100001101010000",  -- ROS word fb2
   "1000000000010000000010000000000000001000011000011111011010000000000011001100000000000010100010001000",  -- ROS word fb3
   "0000000000000000000000000000001011110000000101000001000000000011001110000000000000000100000100000000",  -- ROS word 034
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 035
   "0000000000000111100000000001000000000000000000000111010000000100110110000000001010011001101001001000",  -- ROS word 036
   "1000000000000010000000000000100000000001101000001001001000000000000000000000000000000000101100000000",  -- ROS word 037
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b4
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b5
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b6
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b7
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 134
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 135
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 136
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 137
   "0000000000000110000010000110011000000000000000010011101011111100000010000000000000000100000011100000",  -- ROS word 1b4
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 1b5
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 1b6
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 1b7
   "1000000000000111100010000100110100110000000000000100000101100100000010000000000000000100000100000110",  -- ROS word 234
   "0000000000000111100010000100110100000000000000000100000111100100000010000000000000000000000100000101",  -- ROS word 235
   "1000000000000111100000000000001100010000000000000111000111100100000000000000000000000100000000000100",  -- ROS word 236
   "0000000000000111100000000000001100100000000000000111000111100100000010000000000000000000000000000111",  -- ROS word 237
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2b4
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2b5
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2b6
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2b7
   "1000001001000000000000000001110000000000000000001001001010000100000000000000000000000000000100000000",  -- ROS word 334
   "0000001001000111100010000000110000000000000000001011001010000100000010000000000000000000000100100010",  -- ROS word 335
   "0000000100001100011110000110110000000000000000010010000100000000100101001100100000011010011101110000",  -- ROS word 336
   "1000000100001100011110000110110000000000000000001101011110000000000011001100100000011110011101110000",  -- ROS word 337
   "0000001001000000011110000001110000000000000000001000011000000011001101000100000000000000000100000000",  -- ROS word 3b4
   "1000001001000000000000000001110000000000000000000111000100000100010100000000000000000000000100000000",  -- ROS word 3b5
   "1000000000000000000010000001110101100000000000000111010101101100010010000000000100000000010000100000",  -- ROS word 3b6
   "1000000000000000001010000000000000000000001000000110010100000100000010000000000000000100000100000000",  -- ROS word 3b7
   "1000000000000000000010000000000000000000000000010010011000000001100000000000000000000100000100000000",  -- ROS word 434
   "0000000000000000000010000000000000000000000000001101000101101001100000000000000000000000000100000000",  -- ROS word 435
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 436
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 437
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4b4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4b5
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4b6
   "1000001001000000000010000000000000000000000000010000001010000000000000000000000000000001000000000000",  -- ROS word 4b7
   "0000000000000111100000000000000110100000000101100111011100000100000000000000000000000100110100110000",  -- ROS word 534
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 535
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 536
   "0000000000000111100010000000000000000000000000101001011010000100000010000000000000110101011000000000",  -- ROS word 537
   "1000000000000110000010000000000000000000000101001110011100000100000001011000100000000010110000110000",  -- ROS word 5b4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 5b5
   "0000000000000111000000000000000000000001111000000000001000000000000001011000100000000010000000000000",  -- ROS word 5b6
   "1000000000001001000010000000000000000000000010000000001000000000000000000000000000000100000100000000",  -- ROS word 5b7
   "0000000000000100100000000100110000000000000000110011011000000100000010000000000000000100000100000000",  -- ROS word 634
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 635
   "1000000000000000000000000001000000000000000000001100011010000000000000000000000000000000000100000000",  -- ROS word 636
   "1000000001000111100000000000000000000000000101001010011010000100000010000000000000000000110100110000",  -- ROS word 637
   "0000001010000111100010000000000000000000000000010000011010000000011010000000000000010000010100000000",  -- ROS word 6b4
   "1000000000000000000000000100110000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 6b5
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 6b6
   "0000000000000111100010000000000000000000000101010011011100000100000000000000000000000000110100110000",  -- ROS word 6b7
   "1000000000000010000000000000000000000001111000001101010010110010100000000000000000111001011100000000",  -- ROS word 734
   "0000000000000010000000000000000000000001111000001101010010110000000010000000000000111101011100000000",  -- ROS word 735
   "1000000000010010011000000000000000000011010000101110000110000000000000000000000010000100000000000000",  -- ROS word 736
   "0000000000000000000010000101110000000000000000010010100110000000010010000000000000000000000100110000",  -- ROS word 737
   "0000000000100000001101010000000000000000000000000100000000000011110010000000000000000100000100000000",  -- ROS word 7b4
   "0000001010000000000000000100110000000000000000000000001000000000000000000000000000110000010000000000",  -- ROS word 7b5
   "0000000000000010000010000000000001000011011001001110011010000100000000000000000010000100000000000000",  -- ROS word 7b6
   "1000000000000000000010000110011000000000000000001110011010000100000010000000000100000100000100000010",  -- ROS word 7b7
   "0000000000001010000011100000000000000000000000001111011010000000101000000000000000000000000100000000",  -- ROS word 834
   "0000000000001010000010000000000000000000000000001111011010000000101000000000000000000000000100000011",  -- ROS word 835
   "0000001011000101100010000000000000000000000000010001100000000000000000000000000000000000000100000011",  -- ROS word 836
   "0000000000000010000000000000000000000011011101001111011010000100000010000000000100000000111011100000",  -- ROS word 837
   "0000001010000000100000000000000000000001111110010010011010000000001110000000000000000100110100110000",  -- ROS word 8b4
   "0000001010000000100000000011011000000001111110010011010110000100011010000000000000000100110100110000",  -- ROS word 8b5
   "0000001011010101100010000000000000000011010000010001011000000100000000000000000000000000000100000011",  -- ROS word 8b6
   "0000000000000000000000000101111000000000000101001110011100000000000000000000000000000100000100000000",  -- ROS word 8b7
   "0000000000001010000000000100110010010000000000010001010110000100011110000000000000000100000100000000",  -- ROS word 934
   "0000000000001010100010000100110000000001111000010001010110000100011110000000000000000100110011100000",  -- ROS word 935
   "1000001001000000000010000110110000000000000001010010011100000100000010000000000000000100000100000000",  -- ROS word 936
   "1000000000000111000000000000000000000000000000000110100100000000000001001100000000000100000000000000",  -- ROS word 937
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9b4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9b5
   "1000000000000000000010000000000000000000000000010010010110000100000000000000000000000100000111110000",  -- ROS word 9b6
   "0000000000000010000000000000000000100001011000010011100110100100000000000000000000000100000100000000",  -- ROS word 9b7
   "1000000001000000000000000011101000000000000000010100011010000000010100000000000000111001011100000000",  -- ROS word a34
   "0000000001000000000000000011110000000000000000010100011010000100000000000000000000000100000100110000",  -- ROS word a35
   "0000000001000000000000000000000000000000000000010100011010000100010100000000000000111101011100000000",  -- ROS word a36
   "0011010000100000000000000000000000001000011000010100011000000100000010000000000000000100000100000000",  -- ROS word a37
   "0000001010000000000000000010000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word ab4
   "1000000000010000000000111000000000000011010000010110000111000010100010000000000000000000000100000000",  -- ROS word ab5
   "1000000000001111000000000001110000000000000100110101011010000100000010000000000000000100000001000000",  -- ROS word ab6
   "1000001010000000000010000110000000000000000000110101011100000000000010000000000000010100010100000000",  -- ROS word ab7
   "1000000000000000000010000001001000000000000000010110011000000100000000000000000000000100000100000000",  -- ROS word b34
   "0000000000000010000010000000000001000011011001010110011100000000000010000000000010000100000000000000",  -- ROS word b35
   "1000000000000000000000000001000000000000000000010110011000000101100010000000000000000000000100000000",  -- ROS word b36
   "1000000000010111100010000000000000000011010101010110011100000000000000000000000000000100110100110000",  -- ROS word b37
   "0000000000000000000010000000000000000000000001010111011010000000000010000000000000000000000100000000",  -- ROS word bb4
   "0000000000000000000010000000000000000000000000010111011000000101001000000000000000000000000100000000",  -- ROS word bb5
   "1000000000000111000000000000000000000000000011010111011010000100000011001100000000000010000100000000",  -- ROS word bb6
   "1000000000000000000010000011101000000000000101001000100000000100000010000000000000000100000100000000",  -- ROS word bb7
   "0000100001100000011000010000000010000010001000011000010000000100000001110110110000000111000111010000",  -- ROS word c34
   "1000000001110000011110000110011000000101000000011000011100000000000011110100000000000100110100110000",  -- ROS word c35
   "0000000000000111100000000110111000000000000000011000011010000000000000000000000000000000000000001000",  -- ROS word c36
   "0000001011100000010110010110111000000010001000011000011010000000010100000010000000000000000101000000",  -- ROS word c37
   "1000000000000111000010000100001000001101101000011001011010000000000010111100110000000011001000000000",  -- ROS word cb4
   "1000001011100000011000100110110000000010100000011000100010000000010010000011100001000100000001000000",  -- ROS word cb5
   "0000000001110000000000000000000000000110000000011110011000000100000010000000000000000101011111010000",  -- ROS word cb6
   "0000000000000110000010000110000000000000000000011000101000000000000001001100000000000101000010011000",  -- ROS word cb7
   "0000001011000000000000000000000000001100000000011010011110000100000010000000000000000000000000001000",  -- ROS word d34
   "1000000001100000011100000110011000000110000000011010100010000100000001111100001110000111000011100000",  -- ROS word d35
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d36
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d37
   "1000001010010000011001001110101000000100100000011011101000000110001010000011100001000100000001000000",  -- ROS word db4
   "1000000000000111100000000001000000000000000100111011011010000100000000000000000000000101101000110000",  -- ROS word db5
   "1000001010000000011100110000000000000000000001011011011100000001011010000000100001000100010001001000",  -- ROS word db6
   "0000000000000000000000000111011000000000000011111011011100000100000010000000000000000100000100000000",  -- ROS word db7
   "0000000000001011100000000101101000100000000000011100011010000000000010000000000000010000000000000000",  -- ROS word e34
   "0000000000000010000001010110011000001110010000011111001010000000000010000000000000000100000100000000",  -- ROS word e35
   "0000000000000111100010000101110000000000000101011100010010000110001000000000000000000100000001000000",  -- ROS word e36
   "1000001011001111010101100000000000000000000000011101011111010100000010000010100001110100000000000000",  -- ROS word e37
   "0000000000000010000010000000000000001100100000011001101000010100000000000000000000000001011101000000",  -- ROS word eb4
   "0000000001000000000000000000000000000000000000011110010010000000000000000000000000000101011100100000",  -- ROS word eb5
   "1000000000000111100000001000000000000000000000011000010100000000000000000000000000000100000000100000",  -- ROS word eb6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word eb7
   "0000000000000111100010000110101000000000000000011110011010000100011110000000000000000101101000110000",  -- ROS word f34
   "1000001010000000000010000010111000000000000000011110011000000000011010000000000000000000010001001000",  -- ROS word f35
   "1000000000000000000001010001000000000000000000011111001100010100000000000011110000000000000100000000",  -- ROS word f36
   "0000000000000000000010000000000000000000000101011110011100000000000000000000000000000000000100000000",  -- ROS word f37
   "1000000000100000000000011000000000000110110000011111100000000000000000000000000000000100000001011000",  -- ROS word fb4
   "1000001010010000000001111000000000001000001000011111010110000100000010000011100001000100010001001000",  -- ROS word fb5
   "0010100000000000000010000110110000000000000000011111011010000100000010000000100001000101110011000000",  -- ROS word fb6
   "1011100000001111100010000000000000000000000000011111011100000000000000000000100001000100000100000000",  -- ROS word fb7
   "0000001010000000100010000100110010010001111110000000001100000100011110000000000000000000110100110000",  -- ROS word 038
   "0000000000000000100000000000000000000001111000001101010010110000000010000000000000000100000100000000",  -- ROS word 039
   "0000000000000000000010000000000011110000000000000111001110000000000010000000000000000000000100000000",  -- ROS word 03a
   "0000001101100000000000000000000000000001110000010010011100000100000000000000000000000100101100000000",  -- ROS word 03b
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b8
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0b9
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0ba
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0bb
   "0000000000000000000010000000000000000000000000001110000101111100000000000000000000000000000100000000",  -- ROS word 138
   "0000001011000000000000000110011000000000000000001011011101111100000000000000000000000000000011100000",  -- ROS word 139
   "0000001011000000000000000110011000000000000000001011011101111100000000000000000000000000000011100000",  -- ROS word 13a
   "0000001011000000000000000110011000000000000000001011011101111100000000000000000000000000000011100000",  -- ROS word 13b
   "0000000000000000001010000000000000000001011000010011010011111100000000000000000000000100000011100000",  -- ROS word 1b8
   "1000000000000111111100000000110000000011011000000111100101111100000010011101100000000000000111100000",  -- ROS word 1b9
   "1000000000000111111100000000110000000011011000000111100101111100000010011101100000000000000111100000",  -- ROS word 1ba
   "1000000000000111111100000000110000000011011000000111100101111100000010011101100000000000000111100000",  -- ROS word 1bb
   "0000000000000010000000000000000000000000000101110011100001010100101000000000000000000100000100110011",  -- ROS word 238
   "1000000000000111000010000000000000010000000011001001001000000000000000110000100000000000000000000000",  -- ROS word 239
   "1000000000000011100000000000000000000000000101110011100001010100101000000000000000000100000000110010",  -- ROS word 23a
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 23b
   "1000001010000100111110000101111000000000000100000111001100000100000010000000000000000100000111100001",  -- ROS word 2b8
   "0000001010000100111110000101111000000000000100000100000100000100000010000000000000000000000111100001",  -- ROS word 2b9
   "0000001010000100111110000101111000000000000100000100000100000100000010000000000000000000000111100001",  -- ROS word 2ba
   "0000001010000100111110000101111000000000000100000100000100000100000010000000000000000000000111100001",  -- ROS word 2bb
   "1000000000000000001000000101101000000000000000001011100110000000010000000000000000000000000100000000",  -- ROS word 338
   "0000000000000000001000000101101000000000000000001011100110000000010100000000000000000100000100000000",  -- ROS word 339
   "1000000000000111100000000000000110100000000101101000011100000000000000000000000000000000110100110000",  -- ROS word 33a
   "1000000000000010000000000000100011100000000000000000101000000100000000000000000000001001011101100000",  -- ROS word 33b
   "0000001010000000000000000101111000000000000000001011001110000100010010000000000000000001000000000000",  -- ROS word 3b8
   "1000000000000100100000000110001000000000000101000100011100000000000010000000000000000000000100000000",  -- ROS word 3b9
   "1000000000000000000000000011010110000000000010000110011100000100000000000000000000000000000100000000",  -- ROS word 3ba
   "0000000110100000000010000000000000000001110000000110011100000100000010000000001010000001001100000000",  -- ROS word 3bb
   "1000000000000000000010000001001000000000000010001010011010010100000000000000000000000100000100000000",  -- ROS word 438
   "1000000000000111100000000000010000000000000000001100001000000000000010000000000000000100110000100000",  -- ROS word 439
   "1000000000000000000000000000010000000000000000001100001000000110101000000000000000000000000100000000",  -- ROS word 43a
   "1000000000000000000000000000010000000000000000001100001000000110101000000000000000000000000100000000",  -- ROS word 43b
   "1000000000000110011100000000000110110000000000001011011010000000000000000000000000110101000000000000",  -- ROS word 4b8
   "0000000000000100100000000110001000000000000000110001100000000011001100000000000000000100000100000000",  -- ROS word 4b9
   "0000000000000111111100000000000000000000000000001010011011111100000001001100000000110101000100000000",  -- ROS word 4ba
   "0000000000010010000000000000000011100001100000000000101000000000000000000000000000001101011101100000",  -- ROS word 4bb
   "1000000101000000011100110000110111100000000000001101010110000111110111111101100100000000000100000000",  -- ROS word 538
   "1000000000000110000010000000000000000000000101001101011100000100000001011000100000000010110000110000",  -- ROS word 539
   "1000000110001000100010000000000000000000000000000000001000000000000000000000000000000000000000010000",  -- ROS word 53a
   "0000000000000000000000000000100000000000000000001001001000000000000000000000000000000000000011100000",  -- ROS word 53b
   "1000000000001101000010000111011000000000000000100011000000000011001110000000000000000100000100000000",  -- ROS word 5b8
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 5b9
   "0000000000000000000010000000000000000000000000101100011000010100000000000000000000000000000100000000",  -- ROS word 5ba
   "0000000001100000000000000000000000000001110000001010001110000000000010000000000100000100111101100000",  -- ROS word 5bb
   "1000001001000000001000000110110000000000000000010010011010000100000010000000000000000000000100000000",  -- ROS word 638
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 639
   "1000000000000111000010000110100000000000000000010010011000000101001111001100000000000000000000000000",  -- ROS word 63a
   "0000000000100000000000000000000000000001100000001011011100000100000010000000000000000100000100000000",  -- ROS word 63b
   "1000000000000000000000000110111000000000000000001100011100000000000000000000000000000000000100000000",  -- ROS word 6b8
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 6b9
   "1000000000000000000010000001001110110000000000001011011010010100000000000000000000000100000100000000",  -- ROS word 6ba
   "0000000000000010000000000000000000000001111000001001001000000000000000000000000000000001011000000000",  -- ROS word 6bb
   "0000000000000000000000000011010000000000000011001101011100000000000000000000000100000100010110100000",  -- ROS word 738
   "0000000000000000000000000000000011010000000000000000001000000000000000000000001000000000000000000000",  -- ROS word 739
   "1000000000000000000010000000000110110000000000001010011100000000000010000000000000000100000100000000",  -- ROS word 73a
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 73b
   "0000000001000000000010000101111000000000000000000111011100000000000010000000000000000000000100000011",  -- ROS word 7b8
   "0000000000000000011000000000000011100000000000001110011100000000000010000000000010000000000000000000",  -- ROS word 7b9
   "0000000000000010000010000111011000000000000000001001011101111100000000000000000000000101011000000000",  -- ROS word 7ba
   "0000000000000010000000000000000000000000000000001010001000000000000000000000000000000001000000000000",  -- ROS word 7bb
   "1000000000000111000010000011010000000000000011001011100110000000000011001100000100000000010010100000",  -- ROS word 838
   "0000001010000010000000111000000000000010011000010000011101000000000010000000000000000100000100000000",  -- ROS word 839
   "1000000000000000011110000001000000000000000000110000011000000100000001001110110000000010000000000000",  -- ROS word 83a
   "1000000000000000000010000000000000000000000000010001001000000100000000000000000000000100000100000000",  -- ROS word 83b
   "0000000000000000000000000110001000000000000101010000011100000000000000000000000000000100000100000000",  -- ROS word 8b8
   "1000001010000000000000000011001000000000000000001101010010000000000000000000000000010000010100000000",  -- ROS word 8b9
   "0000001001000100100010011000000000000000000001010000011100000100000000000000000000000101000000000000",  -- ROS word 8ba
   "0000001011100000000010000000000000000001100000001101100100000100000010000000000000000000101100000000",  -- ROS word 8bb
   "0000000000000000011100000000000000000000000000001001001000000000000000010100100000000000000000000000",  -- ROS word 938
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 939
   "1000000110010000000000000000000000000001100000000101100110000100000010000000000000001001001111100000",  -- ROS word 93a
   "1000000000000111000000000000000000000000000000010011011000000100000001001100000000000100000000000000",  -- ROS word 93b
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9b8
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9b9
   "1000000000000100100000000101001000000000000001001101100100000000000010000000000000000000000100000000",  -- ROS word 9ba
   "1000000000100000000011010000000010010000100000010011011111000000000000000000000000000100000100000000",  -- ROS word 9bb
   "1000000000000000000010000000000000000001111000010100011100000100010100000000000000000100000100000000",  -- ROS word a38
   "0000000001000000000000000000000000000000000000010100011110000000000000000000100000000100000101000000",  -- ROS word a39
   "1000000000100000000111010100010000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word a3a
   "0000000000100000000101010100000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word a3b
   "1000000000000000000010000000000000000000000011110110001000000010100010000000000000000100000100000000",  -- ROS word ab8
   "0000000001000000000000000000000000000000000000010101011100000100000010000000000000000100010100100000",  -- ROS word ab9
   "0000001010000000000010000000000000000000000011110101001010000000000000000000000000000100000000001000",  -- ROS word aba
   "1000000000000100100010000000011000000011011000010100100110000100010100000000000000000101011111010000",  -- ROS word abb
   "1000000000000010000000000000000000000000000000010110011010010100000000000000000000000100000000001000",  -- ROS word b38
   "0000000000010010011000000000000000000011010000110110100010000000000010000000000010000000000000000000",  -- ROS word b39
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b3a
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b3b
   "0000000000000010000010000111101000000000000000010110001100000100000010000000001010000000000100110000",  -- ROS word bb8
   "0000000000000010000000000000101000000000011000110110010000000100000000000000000000000100000100000000",  -- ROS word bb9
   "0000000000000010011100000110110000000000001000010111011100010100000010000011111110000100000100000001",  -- ROS word bba
   "0000000000000010000000000000000000000000000000110110010000000100000000000000000000000100000100000000",  -- ROS word bbb
   "1000000000000010000000000000000000001101100000011001000110000001100100000000000000000101000000000000",  -- ROS word c38
   "0000000000000111100010000000101000000000000000011000011110000100000001010000110000000010000111100000",  -- ROS word c39
   "0000000000010111100000000110011000010101010000111000011000001110100010000010110000000100000100001000",  -- ROS word c3a
   "1000000000010111100000000100101000000101010000111001001000001100000010000000000000000100110000001000",  -- ROS word c3b
   "1000000000000110000010000110000000000000000000011000101000000000000001001100000000000101000110001000",  -- ROS word cb8
   "1000000000000110011100110001111000000000000000011000011110100000000011001000100001000100000000001000",  -- ROS word cb9
   "1000000001010000000000000000000000000110100000011001001010000010100010000000000000000100000001000000",  -- ROS word cba
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word cbb
   "0000001010000000000010000110110000000000000011011011011010000000000010000000000000000100010001001000",  -- ROS word d38
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d39
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d3a
   "1000000000010010000000000000000000000100000000011010011110000000000010000000000000000101000000000000",  -- ROS word d3b
   "1001010000001011100010000000000000000000000000011011010010000100000010000000000000000100000100000000",  -- ROS word db8
   "0001010000101011100000000110011000000101011101011011011010000100000010000000000000111000000000000000",  -- ROS word db9
   "1000000001000010000000010000000000000000000000011010000000000110001000000000000000110101011000000000",  -- ROS word dba
   "0000000000000110000001100000000000001101011000011011010010000100000010000010100001000100000111100000",  -- ROS word dbb
   "1001010000001010000010000100111000000000000000011100011010000000000000000000000000000100000100000000",  -- ROS word e38
   "1000000000011111000010000110011000000011010000011101010010000000000000000000000000000100000100000000",  -- ROS word e39
   "0000000000000111100010000001001000000000000100111100100100000100000010000000000000000000110100110000",  -- ROS word e3a
   "1000000000010000000000000000000000000100100000011100100100000000000000000000000000000000000100011000",  -- ROS word e3b
   "1000001011000011000011100000000000001101011000011110001010000100000000000000100001000000000011100000",  -- ROS word eb8
   "0000000000000011000001100000000000001101011000011101100110000100000010000000100001000000000011100000",  -- ROS word eb9
   "0000000000000010000000000000000000001100101000011100000100000100000010000000000000000100000100110000",  -- ROS word eba
   "1000000000000000000010011000000000000000000000011101011100000110001000000010001000000100000100101000",  -- ROS word ebb
   "0000001001000000000001010001000000000000000001011111001100010100000000000011110000000100000100000000",  -- ROS word f38
   "1000000001010000000000000111011000000100111000011110011110000010001001001100000000000110000000001000",  -- ROS word f39
   "1000000000000010000000011001111000001100000000111110011100000000000011010000100001000010001100000000",  -- ROS word f3a
   "0000000000000010010110110110011000001100001000111101010010000100000000000000100001000100000000001000",  -- ROS word f3b
   "0010110000100000011111010000000000001000000000011111011010000001101110000000001010000001001100110000",  -- ROS word fb8
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fb9
   "0000000000000000000010000000000000000000000000011111010010011000000000000000000000000000000100000000",  -- ROS word fba
   "0000000000000000000010000000000000000000000100111111010110000000000010000000000000000000000100000000",  -- ROS word fbb
   "0000000110000000000010000000000000000000000000001010001001001100000000000000000100000100111001000000",  -- ROS word 03c
   "1000000000000000000010000000000000000000000000010001010100110000000000000000000000000101011111010000",  -- ROS word 03d
   "1000000000010000000010000000000000000011010000001101000110000100000000000000000000000100000100000000",  -- ROS word 03e
   "0000000000001001000010000000000000000000000000010011000110000000000000000000000000000000000100000000",  -- ROS word 03f
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0bc
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0bd
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0be
   "1000000000000000000000000010011000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 0bf
   "0000001011000000000000000000000000000000000000001000010101111100000010000000000000000000000011100000",  -- ROS word 13c
   "0000001011000000000000000110011000000000000000001011011101111100000000000000000000000000000011100000",  -- ROS word 13d
   "0000001011000000000000000110011000000000000000001011011101111100000000000000000000000000000011100000",  -- ROS word 13e
   "0000001011000000000000000110011000000000000000001011011101111100000000000000000000000000000011100000",  -- ROS word 13f
   "1000000000000111111100000000110000000000000000000011100111111100000011111101100000000000000111100000",  -- ROS word 1bc
   "1000000000000111111100000000110000000000000000000001100101111100000010011101100000000000000111100000",  -- ROS word 1bd
   "1000000000000111111100000000110000000011011000000111100101111100000010011101100000000000000111100000",  -- ROS word 1be
   "1000000000000111111100000000110000000011011000000111100101111100000010011101100000000000000111100000",  -- ROS word 1bf
   "1000000000000010000000000000000000000000000101100100011110000000000010000000000000000000000100110011",  -- ROS word 23c
   "1000000000010000000000000000000011110000101000000111001000000100000010000000000100000100010011010000",  -- ROS word 23d
   "0000000000000011100000000000000000000000000101100100011110000000000010000000000000000000000000110010",  -- ROS word 23e
   "0100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 23f
   "0000001010000100100000000101111000000000000100000100000010000100000000000000000000000100000111100001",  -- ROS word 2bc
   "0000001010000100100000000101111000000000000100000100000010000100000000000000000000000100000111100001",  -- ROS word 2bd
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2be
   "0000000000100000000000000010011000000011010000000111001100000000000010000000000000000100000100000000",  -- ROS word 2bf
   "1000000110000000001000000000000000000000000000000000011010000100000010000000000100000000111101100000",  -- ROS word 33c
   "0000000000000000011100000000000000000000000000001011100100000011001010000011100000000000000000000000",  -- ROS word 33d
   "1000000000010010000010000110111000001011110000010111001000000000000000000000000000111000000000000000",  -- ROS word 33e
   "1000000000000000000000000101001000000000000000010000001110000100000000000000000000000000000100000000",  -- ROS word 33f
   "0000000000100000000000000000000000000001100000000110011110000000000000000000000000000100000100000000",  -- ROS word 3bc
   "1000000000000010000000000000000000000001111000001010001000000000000010000000000000000100000011010000",  -- ROS word 3bd
   "0000000000000111000010000110100000000000000101001111100100000100000011001100000000000100000000000000",  -- ROS word 3be
   "1000000000000010000010000000000000000001011000010011010010000000000000000000000000000000000001000000",  -- ROS word 3bf
   "0000000001000000000010110000100000000000000000001010001110000000100000000000000100000101111000000000",  -- ROS word 43c
   "1000000000010010111100000110011000000011010000001011100010000000000010000000100000000100101011110000",  -- ROS word 43d
   "0000000000000000000000000110001000000000000011000111011110000100000000000000000000000100000100000000",  -- ROS word 43e
   "1000000000000010100000000000000000100001001000010010010010000000000000000000000000000101010001000000",  -- ROS word 43f
   "0000000001000000000010110000100000000000000000001010001110000000100000000000000100000100111001000000",  -- ROS word 4bc
   "1000000000000010111100000110110000000000000000001011100010000000000010000000100000000100101011110000",  -- ROS word 4bd
   "0000000000000000000000000110001000000000000101001111100100000100000010000000000000000100000100000000",  -- ROS word 4be
   "0000000000000010000000000000000000000001111000001011100110000000000010000000000000000001011000000000",  -- ROS word 4bf
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 53c
   "1000000000000010111100000000000000000000000000010010000110000100000010000011100000000100000000000000",  -- ROS word 53d
   "0000000000000111000000000000000000000001111000001011100110000000000011001100000000000000000000000000",  -- ROS word 53e
   "0000000110000111000010010110110101000000000000001100000000000100000011001100000000001110101000000000",  -- ROS word 53f
   "1000000101000000000010110000000111100000000000001011010010000011110110000000000100000000000000000000",  -- ROS word 5bc
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 5bd
   "1000001001000000001000000000000000000000000000001010011110000100000000000000000000000000000100000000",  -- ROS word 5be
   "0000000000000000000010000000000000000000000000010000100110000100000110000000000000000000000100000000",  -- ROS word 5bf
   "1000000000000010111100110000110111100000000000001011011110000000000001111101100000000001110100000000",  -- ROS word 63c
   "1000000100001100011110000000000000000000000000001111100010000100000011001100100000011110011101110000",  -- ROS word 63d
   "0000000000000000000000000110010000000000000000001011011110000100000000000000000000000100000100000000",  -- ROS word 63e
   "0000000000000000000010000000000000000000000000001011011110000100000010000000000000000000000100000000",  -- ROS word 63f
   "1000000000000111111100000000110000000000000000000011100100000000000011111101100000000000000101000000",  -- ROS word 6bc
   "1000000100001100011110000001111000000000000000001100011110000000000010111100100000011010011001110000",  -- ROS word 6bd
   "0000000101001100000000000110001000000000000000001111000010000100101100000011100000000000101000000000",  -- ROS word 6be
   "1000000000000010000000000000000000000000000000001100011110000100000010000000000000000100000011010000",  -- ROS word 6bf
   "0000000000001101001010000000000000000000000000010010100000000011001100000000000000000000000100000000",  -- ROS word 73c
   "1000000000010010000000000000000000000011010010001011100110000000000010000000000000000101011000000000",  -- ROS word 73d
   "1000000101000000011110000110101101010000000000010011100100000000000010000000000000000101100111000000",  -- ROS word 73e
   "0000001011001101000010000000000000000000000000001101000010000101001100000000001010000101000000000000",  -- ROS word 73f
   "1000000000000000000000000101010000000000000000010000010101010100000010000000000000000000000100000000",  -- ROS word 7bc
   "1000000000000010000000000000000000000011011101001110011110000000000010000000000000000101000000000000",  -- ROS word 7bd
   "1000000101000000011110000110101101010000000000010011100100000000000010000000000000000101100111110000",  -- ROS word 7be
   "0000000000001100001000000000000000000001111000001001000100000100101101001101010000000010001000000000",  -- ROS word 7bf
   "1000000000000000000010000110101000000000000000001100011000001100000011001010000000000000000000000000",  -- ROS word 83c
   "1000000100000000000000000000000000000000000000001111011110000000000010000000001010000001100100000000",  -- ROS word 83d
   "1000000101000000011110000110101101010000000000010011100100000000000010000000000000000101100100000000",  -- ROS word 83e
   "1000000110000000011100110000000000000000000000001111011110000100000011001101010100001110001000000000",  -- ROS word 83f
   "0000000000100000001100000000000000000000000000000100000000000011110010000000000000000100000100000000",  -- ROS word 8bc
   "0000000100001100011110000110101000000000000000001111100010000110000011001100100000011010011101110000",  -- ROS word 8bd
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 8be
   "0000000000000000001000000000000000000001111000001001001010000000000110000000000000000100000100000000",  -- ROS word 8bf
   "0000000000000010000000000011011000000001111000010011101010000100011110000000000000110001011000000000",  -- ROS word 93c
   "0000000100001100011110000000000000000000000000001111100010000100000011001100100000011110011000000000",  -- ROS word 93d
   "0000001101000010100000000000000000000000000000010011101010000000000000000000000000000100101100000000",  -- ROS word 93e
   "1000000000000000001000000000000000000001111000001001001000000000000110000000000000000000000100000000",  -- ROS word 93f
   "0000000000000000000010000000000000000000000000000000001001100000000000000000000000000000000100000000",  -- ROS word 9bc
   "0000000000000000000000000000000110100000000101110011011110000100000010000000000000000100000100000000",  -- ROS word 9bd
   "1000000000000000000010000000000000000000000000000000001000000011001110000000000000000100000100000000",  -- ROS word 9be
   "1000000000000000000010000000000000000000000010001001100011010100000000000000000000000100000100000000",  -- ROS word 9bf
   "1000000000000010000000000000000000000000000000010100011110000110001000000000000000000000000100000000",  -- ROS word a3c
   "1001000000000000011100000110100000000000000000010100100000000000101110111100000000000000000100000000",  -- ROS word a3d
   "1000000000000000011100000000000000000011011000010100011110000000000011000100000000000000000100000000",  -- ROS word a3e
   "0000000000100000000101010100011000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word a3f
   "1000000000000010000000000110101000000000000000010101011110000100000011001000100000111000110100000000",  -- ROS word abc
   "0000000000000010000010000110010000000000000000010101011111111100000000000000000000000100001000000000",  -- ROS word abd
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word abe
   "0000000000010010000010000110101000000001100000010100010000000010001001001000100000011010000100000000",  -- ROS word abf
   "0000000000000000000000111000000000000000000000010110011000000000000010000000000000000100000100000000",  -- ROS word b3c
   "1000000000000111100010000101101000000000000000010110100000000011011000000000000000000100110100110000",  -- ROS word b3d
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word b3e
   "0010000000010111100010000000000010001000000000010111100000100000000010000000000000000000110100110000",  -- ROS word b3f
   "1000000000000000000010000000000000000000000000010111011000000001001000000000000000000100000100000000",  -- ROS word bbc
   "0000000000000100100010000000000000000000000000110111100110011000000010000000000000000000000100000000",  -- ROS word bbd
   "0000000000000000000010000000000000000000000000010111100100011100010100000000000000000000000100000000",  -- ROS word bbe
   "1000000000100000000111010011110000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word bbf
   "0000000000000010000010000000000010001101001000011001000110000100000000000000000000110101011000000000",  -- ROS word c3c
   "1000001011000000000000000110000000000000000000011001001010000100000000000010001010000100000001100000",  -- ROS word c3d
   "0000000000000010000010000000000000001101000101011001000000000100000010000000000000000000000100110000",  -- ROS word c3e
   "1000001011000000000000110110000000000000000000011001001010000110001001010000101011000110000001100000",  -- ROS word c3f
   "1000001011000010000000011110101000001101101000011001011000000010001001010011100001000010000110011000",  -- ROS word cbc
   "0000000000000000000000000001000001010000000000011001100000000000001100000000000000000100000100000000",  -- ROS word cbd
   "0000000000000010011000011001111000000000000000011010100100000100000010000011100001000000000010011000",  -- ROS word cbe
   "0000000000000000000010000000000000000000000000011001100100000100011010000000000000000000000100000000",  -- ROS word cbf
   "0011110000000010000000000000000000001100101000011010010010000100000000000000000000000101011100111000",  -- ROS word d3c
   "0000000000000000011101010101101000001100000000011010011110000100000000000011100001000100000100000000",  -- ROS word d3d
   "0000001011010000011100000000000000000100001000011010100100000000000001111100000000000010000001000000",  -- ROS word d3e
   "0000000000000010000010000000000000001100001000011010000110000100000000000000000000000101011000000000",  -- ROS word d3f
   "0000000000000111000000000000000000000000000000011011011110000000000011010000100000000000000000000000",  -- ROS word dbc
   "0000000000000111011110000000000000000000000000011011011110000100000001001000100000000010000100000000",  -- ROS word dbd
   "0000000000000000011100000000000000000000000000011011011110000100000010011100000000000110000100000000",  -- ROS word dbe
   "1000000000000000011100000000000000000000000000011011100000000100000100011111110000000010000100000000",  -- ROS word dbf
   "0000000000010010000000000000000000001100100000011100100100000000000000000000000000000000010000011000",  -- ROS word e3c
   "0000000000000111100010000000000000000000000100111100100100000100000010000000000000000000110100110000",  -- ROS word e3d
   "0000000000010000000000000001000000000100110000011100100100000100000000000000000000000100000100011000",  -- ROS word e3e
   "0100000000000010000010000000000000001100010000011101010100000100000010000000000000000100010000000000",  -- ROS word e3f
   "1000000000000000000010000000000000001100110000011100001100000000000010000000000000000100000100000000",  -- ROS word ebc
   "0000000000000000010110011101101000001100110000011001101000000000000001000110110000000010000100000000",  -- ROS word ebd
   "0000000000000111100010000000000000000000000000011100011010000100000010000000000000000101011000000000",  -- ROS word ebe
   "1000000000000010000010000000000010001100101000011101010010000100000010000000000000000100000100110000",  -- ROS word ebf
   "1000000000000010000010000110100000000000000000011110011110000110001000000000000000000000010000000000",  -- ROS word f3c
   "1000000000000010000010000000000000001100001000011111000000000000000000000000000000000000001000000000",  -- ROS word f3d
   "1000000000000000011100000100011010000000000000011101010110000000000000000000000000000000000100000000",  -- ROS word f3e
   "0000001010010000000010000110100000000101000000011110010110000000000010000000000000000100000001000000",  -- ROS word f3f
   "1000000000000000000010000000000000000000000000011111011100000101001100000000000000000100000100000000",  -- ROS word fbc
   "0000000000110101100010000000000000000011010000011111011110000010001000000011110000000000000100000000",  -- ROS word fbd
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fbe
   "0000000000010000011100111000000000000010111000011111100000000010001001001111110000000110000100000000",  -- ROS word fbf
   "1000001101000010111110000000000000000000000000000000100000110100101101001111110100000010000011110000",  -- ROS word 040
   "1000000000000010111100000000000000000000000000000000100000110100101101001111110100000010000110110000",  -- ROS word 041
   "0000000101000010111110000000000000100000000000010011100010000011010011111100001100000001110111000000",  -- ROS word 042
   "0000000101000010111110000001001000100000000000001000100010000011010011111100000000000001110111000000",  -- ROS word 043
   "1000000101000000000010000110011000000000000000000111100010000100000010000000000000000001110011000000",  -- ROS word 0c0
   "1000000000000010100010000110011000000000000000000001100100000100000000000000000000000100000111110000",  -- ROS word 0c1
   "0000000100000000011110000110011000000000000000000001100010000100000001001111111010000111110000000000",  -- ROS word 0c2
   "1000000000000010100010000110011000000000000000000001100100000100000000000000000000000100000111110000",  -- ROS word 0c3
   "1000000000010010000010000000000000000001010000000010100000000000000010000000000000000001000000000000",  -- ROS word 140
   "1000000101000000000000000000000000000001011000000010100010000100101100000000000000000000000100000000",  -- ROS word 141
   "0000000100000010011100000001011000000001011000000010100000000011011111001110111010000111110100000000",  -- ROS word 142
   "0000000000000010001010000000000000000001001000010011010010000100000010000000000000000000000100000000",  -- ROS word 143
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 1c0
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 1c1
   "0000000000000010001000000000000000100001001000001111000110000000000000000000000000000100000100000000",  -- ROS word 1c2
   "0000000000010111100000000000000110010011010101001001000000000000000000000000000000000100000100000000",  -- ROS word 1c3
   "1000000000000011000000000101000000000001011000010010010010000000111001001100000000000010000100110000",  -- ROS word 240
   "0000000000000000000010000101000000100001011000010010010010000000000000000000000000000100000010110000",  -- ROS word 241
   "1000000100000010111110000000000000000000000000001000100100000000000001001110111010000011001011110000",  -- ROS word 242
   "0000000000000000001000000001000000000001011000010011100110100100000000000000000000000100000100000000",  -- ROS word 243
   "0000000000000010000000110010110011100001111000000101100100000100100000000000001010001100000111100000",  -- ROS word 2c0
   "1000000000000010000000110010110011100001111000000101100100000100100000000000001010001100000001100000",  -- ROS word 2c1
   "0000000000000010000000110010110011100001111000000101100100000100100000000000001010000100101100000000",  -- ROS word 2c2
   "0000000110000000000000110000000011100000000000000101100100000000100000000000001010001000000001100000",  -- ROS word 2c3
   "0000000000000010000000110000011000000001111000000110100100000000100000000000000100001000000011100000",  -- ROS word 340
   "1000000110000000000010000000000000000000000000000110100110000000000010000000000100001100000101100000",  -- ROS word 341
   "1000000000000010000000000000000000000000000000000110100100000100100000000000000100000100101000000000",  -- ROS word 342
   "1000000000000010000000000000000000000000000000000110100100000000000010000000000100001000000101100000",  -- ROS word 343
   "0000000101000010111110000000000000100000000000001000100100000011010011111100000000000001110100000000",  -- ROS word 3c0
   "0000000000000000001000000000000000000001001000000111011110000100000010000000000000000000000011100000",  -- ROS word 3c1
   "1000001101000010111110000000000000000000000000000000100000110100101101001111110100000010000011110000",  -- ROS word 3c2
   "0000000000001001000000000000000110010000000101000101100110000000000010000000000000000100000100000000",  -- ROS word 3c3
   "0000000000000010111100000001010000000001001000000100100000000011011011001111110100000011100000000000",  -- ROS word 440
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 441
   "0000000000000010111100000001010000000001001000001000100110000111011111001111110100000011100000000000",  -- ROS word 442
   "0000000000000000000010000011110000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 443
   "1000000000000111000010100110000000000000000011001001100100000011000101010100000000000000000000000000",  -- ROS word 4c0
   "0000000000000111000000000000000000000000000000001011100110000110001111010100000000000000000000000000",  -- ROS word 4c1
   "1000000000000000000000000000000010000000000101101100101000010000000010000000000000000000000100000000",  -- ROS word 4c2
   "1000000000000000000000000000000010000000000101101101001000010000001110000000000000000000000100000000",  -- ROS word 4c3
   "0000001010000000000010000000000000000000000100010001001100000000000010000000000000110100010000000000",  -- ROS word 540
   "1000000000000111000010100110000000000000000011001010100000000011000101110000100000000100000100000000",  -- ROS word 541
   "0000000000000000000010000000000000000000000101101001011000010000000010000000000000000000000100000000",  -- ROS word 542
   "1000000000000000000010000000000000000000000101100111011000010000000010000000000000000100000100000000",  -- ROS word 543
   "1000000000000010111100000001001000000000000000001011100010000100000000000011100000000100101011110000",  -- ROS word 5c0
   "1000000000000010111100000000000000000000000000010010000110000100000010000011100000000100101011110000",  -- ROS word 5c1
   "0000000000000010100010000000000000000000000000000110011110000000000011101000000000000010101111110000",  -- ROS word 5c2
   "1000000000000010111100000000000000000000000000010010000110000100000010000011100000000100101011110000",  -- ROS word 5c3
   "0000001101000010000010000000011000000001111000001001011110000000000000000000000100001100000011100000",  -- ROS word 640
   "0000000110000000000010000000000000000000000000010001011100000100000010000000000100001000000101100000",  -- ROS word 641
   "0000000110000000000010000000000000000000000000001100100110000100000000000000000100001100000011100000",  -- ROS word 642
   "1000000110000010000000000000000000000001111000001100011100000100000010000000000100001000000101100000",  -- ROS word 643
   "1000001100100000000010000000000000000001110000000000101000000000000010000000001010000000000011100000",  -- ROS word 6c0
   "1000001000000010000000000000000000000001101000001101100110000100000000000000000000000000000101100000",  -- ROS word 6c1
   "1000000110000000000010000000000000000000000000001101100100000000000000000000000000000000000011100000",  -- ROS word 6c2
   "0000000110000000000010000000000000000000000000000101100110000000000000000000000000000000000101100000",  -- ROS word 6c3
   "0000000000000010000000000000000000000001111000001110100010010100000010000000000000000101011111100000",  -- ROS word 740
   "1000000000000010000000000000000000000001111000001110100010010100000010000000000000000101011000000000",  -- ROS word 741
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 742
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 743
   "0000001011000000000000000000000000000000000000001111100000000100000010000000001010000001000000000000",  -- ROS word 7c0
   "1000000000001101000000000000000000000001111000001011100110000000000010000000000000000000000100000000",  -- ROS word 7c1
   "1000000000000010000010000101100000000000000000001011011000000100000000000000000000000100000100110000",  -- ROS word 7c2
   "0000001011001101001000000000000000000000000000001111100010000001001100000000001010000001000000000000",  -- ROS word 7c3
   "0000000000001001100010000000001000000000000000001100100110000100000010000000000000000000000100000000",  -- ROS word 840
   "0000000000000000000010000000000000000000000000000011101000000100000000000000000000000000000100000000",  -- ROS word 841
   "1000001011000000011010000000000011100000000000001110000000000100000010000000000010000000000000000000",  -- ROS word 842
   "0000000001000000011000000011100011100000000000000011101000000100000000000000000010000000000000000000",  -- ROS word 843
   "1000000000000000011100011000000000000000000000010001100000000100001010000010110000000100000000110000",  -- ROS word 8c0
   "0000000000000111001000000000000000010000000000010010011100000000000001001000100000000000000000000000",  -- ROS word 8c1
   "0000000000000000000000000000000110010000000101010001011100000100000000000000000000000100000100000000",  -- ROS word 8c2
   "0000000000100000000000011000000000000010111000010000011100000100000000000000000000000001000000000000",  -- ROS word 8c3
   "0000000000001101000000000000000000000000000000100011001000000011001100000000000000000100000100000000",  -- ROS word 940
   "0000000101001001000010011000000011000000000000001111100110000000001010000000000000000000000100000000",  -- ROS word 941
   "1000001001000100100010000000000000000000000001001001100011010100000000000000000000000101011101000000",  -- ROS word 942
   "0000000000000000011100000000000000000000000010010011011110000000000010111100000000000010000000000000",  -- ROS word 943
   "0000000000010000000010000000000011110000100000000111000110000100000000000000000100000100010011010000",  -- ROS word 9c0
   "1000000000010000000010000000000011110000100000000111000110000100000010000000000100000000010011010000",  -- ROS word 9c1
   "1000001010000000000010000000000000000000000000100000001000000000000000000000000000010100010100000000",  -- ROS word 9c2
   "1000000000000000000010000000000000000000000000100000001000000000000000000000000000000100000100000000",  -- ROS word 9c3
   "0001000000000000011110000110110000000000000000010100011110000000000011000100000000000000000100000000",  -- ROS word a40
   "0000000000010000000010000110111000100011010000010101000000000000000000000000000000000000000100000000",  -- ROS word a41
   "0001000000000000011100000110100000000000000000010101000000000000000010111100000000000100000100000000",  -- ROS word a42
   "1000000000000000000010000001111000000000000000010101000000000100000000000000000000000100000100000000",  -- ROS word a43
   "0000000001000000011100000110011000000000001000010101011110000000000010000000100000000100100100000000",  -- ROS word ac0
   "0000000000000000000010000000000000000000000000010101001110000100000000000000000000000000000100000000",  -- ROS word ac1
   "1000000000000000000010000011101000000000011001010100100110000000000000000000000000000100000100000000",  -- ROS word ac2
   "0000000000000000000010000000000010100000000000010101010000000000000010000000000000000000000100000000",  -- ROS word ac3
   "0000000000010000000000000000000010001011101000010111100000000000000010000000000000000100000100000000",  -- ROS word b40
   "0000000000010000000000000001001000001000001000010111100000000000000010000000000000000100000100000000",  -- ROS word b41
   "0011010000010000000000000000000010001010101000010111100000000000000010000000000000000100000100000000",  -- ROS word b42
   "1000000000010000000010011001000000001011111000010111100000000000000010000000000000000100000100000000",  -- ROS word b43
   "0000000000000000000000111000000000000000000010010110000101000000000000000000000000000100000100000000",  -- ROS word bc0
   "1000000000000000000000000101001000000000000000010110011010000000000010000000000000000000000100000000",  -- ROS word bc1
   "1000001010000000000010000000000000000000000010110101001010000000000000000000000000000000000000001000",  -- ROS word bc2
   "1011010000010000000010000101101001011011100000010111100000000000000010000000000000000100000100000000",  -- ROS word bc3
   "0000000000000111100010000000000000000000000000011000100000000100000000000000000000000100000000001000",  -- ROS word c40
   "0000000000000111111100000000000000000000000000011000101010000100000000000000100000000100000100001000",  -- ROS word c41
   "1000001011010000011100000110010000000101010000011000100100000100000000000000100000000001011100000000",  -- ROS word c42
   "0000000000100000010100010110111000000010001000011000011010000000000000000010000000000000000000000000",  -- ROS word c43
   "0000000000000010000000000000000000000000000000011000010110000100000000000000000000000100000101001000",  -- ROS word cc0
   "1000000000000111100010000011100110010000000101011001100000000100000000000000001010011001101001001000",  -- ROS word cc1
   "1000001001000000011100000100111000000000000001011001100000000100000010000000000000000000000100000000",  -- ROS word cc2
   "0000000000000010000010000101101110010011011101111001100010000000000000000000000000101101000000000000",  -- ROS word cc3
   "0000110000000000000010000110110000000000000000011010100010000100000010000000000000000001011111010000",  -- ROS word d40
   "0000001011100000000000000000000000000100000000011010100100000000000000000000000000000001011000000000",  -- ROS word d41
   "0000110000100000000010000110110000000100110000011010100010000010001000000000000000000001011111010000",  -- ROS word d42
   "0000000000000111000010000111011000000000000000011011011110000000000000000010110000000100000000000000",  -- ROS word d43
   "0000001011000000000010010110111000001110011000011011011100000100000001001000110000000101101001001000",  -- ROS word dc0
   "0000000001000000000000000000000000000000000000011010000110000100000010000000000000011001011000000000",  -- ROS word dc1
   "0000000000000000000010000000000000000000000000011011100010000000000001001000100000000100000000000000",  -- ROS word dc2
   "0000001011000111000010000000000000000000000000011011100010000100000011001111110000000110000001000000",  -- ROS word dc3
   "0000000000000010000000000001000000001100100000011100100100000011111010000000000000000000010000011000",  -- ROS word e40
   "1000000000100000000000110000000000000100100000011100100010000011111010000000000000010001011100000000",  -- ROS word e41
   "0000000000000010000010000000000000001100100000011100100100000100000000000000000000000100010000011000",  -- ROS word e42
   "1000000001000000011000000110111000001110000100011100100010000100000010000000000000000100000000001000",  -- ROS word e43
   "1010100000000000000010000110101000000000000000011101101010000110001001010000100001000100000100000000",  -- ROS word ec0
   "0000000000000000000010000001111000000000000101011101101010000000000000000000000000000000000100000000",  -- ROS word ec1
   "0000000000000000010100100110101000000000000000011101100000000000001111010000100001000100000100000000",  -- ROS word ec2
   "1000001010010000000010000010111000000100011011011101100010000000011010000000000000000000010001001000",  -- ROS word ec3
   "1000000000001111000010000000000000000000000000011110101000000100000000000000000000000000000000001011",  -- ROS word f40
   "1000001010000000000010000010111000000000000000011110100010000000011010000000000000000000010001001000",  -- ROS word f41
   "1000000000001111000010000000000000000000000000011110101000000100000000000000000000000000000000001011",  -- ROS word f42
   "0000000000000111100010000110101000000000000000011110011010000100011110000000000000000101101000110000",  -- ROS word f43
   "0000000000000000000010010000000000000010011000011111011110000100000011010010100001000010000100000000",  -- ROS word fc0
   "0011100000000000000000000000000000000000000000011111010100000100000000000000100001110100000100000011",  -- ROS word fc1
   "1000000000000010000010000000000000101100101000011100011000000000000010000000000000000101000111100000",  -- ROS word fc2
   "0000000000000010000000000001000000101100101000011100011000000000000010000000000000000101000111100000",  -- ROS word fc3
   "0000001101000010111110000000000000000000000000000000100010110100101101001111110100000110000011110000",  -- ROS word 044
   "0000000000000010111100000000000000000000000000000000100010110100101101001111110100000110000110110000",  -- ROS word 045
   "1000000101000010111110000000000000100000000000001000100000000011010011111100000000000101110111110000",  -- ROS word 046
   "1000000101000010111110000001001000100000000000001000100000000011010011111100000000000101110111110000",  -- ROS word 047
   "1000000101000000000010000000000000000000000000000111100010000100000010000000000000000001110011000000",  -- ROS word 0c4
   "1000000001100000011110000001111000000010000000000001100000000011110111001110000000000110000111100000",  -- ROS word 0c5
   "0000000100000000011100000001011000000000000000000001100010000011011111001111111010000011110000000000",  -- ROS word 0c6
   "0000000000000010001010000000000000000001001000010011010010000100000010000000000000000000000100000000",  -- ROS word 0c7
   "1000000100000010011100000000000000000000000000000010100000000100000001001110111010000011110100000000",  -- ROS word 144
   "1000000100000000011110000000000000000000000000000010100000000100000001001110111010000011010000000000",  -- ROS word 145
   "0000000000100000011100110000000111100011010000000010100100000000000001001110000000000010000000000000",  -- ROS word 146
   "1000000000010010000010000000000000000001010000000011100010000000000000000000000000000100000100000000",  -- ROS word 147
   "1000000101000000011100110000000111100000000000000010100100000000101101001110000000000110000000000000",  -- ROS word 1c4
   "1000000000000010100010000000000000000000000000000011100110000100000000000000000000000100000111110000",  -- ROS word 1c5
   "1000000001000000000000000000000000000011011000000010100010000000101100000000000000000100000001000000",  -- ROS word 1c6
   "0000000000000010100010000000000000000000000000000011100100000100000000000000000000000000000111110000",  -- ROS word 1c7
   "1000000000000011000000000101000000000001011000010010010010000000111001001100000000000010000100110000",  -- ROS word 244
   "0000000000000000001010000101000000000001011000001000011110000100000010000000000000000000000100000000",  -- ROS word 245
   "1000001110000010011100000000000000000000000000001000010100000100000001001110111010000111001011110000",  -- ROS word 246
   "1000000000000000000010000001000000000001011000010011100110100100000000000000000000000100000100000000",  -- ROS word 247
   "0000000000000000001000000000011000000000000000000101100100000100000000000000000000000000000011100000",  -- ROS word 2c4
   "1000000000000010001010000010110011100001111000000101100100000100000000000000000000001000000001100000",  -- ROS word 2c5
   "0000000000000010001010000010110011100001111000000101100100000100000000000000000000000000101100000000",  -- ROS word 2c6
   "0000000110000000000000000000000011100000000000000101100010000100000000000000000000001000000001100000",  -- ROS word 2c7
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 344
   "1000000110000000001000000000000000000000000000000110100110000000000000000000000100001000000101100000",  -- ROS word 345
   "0000000000000010001010000000011000000001111000000110100100000000000000000000000100000100101000000000",  -- ROS word 346
   "1000000000000010001010000000011000000001111000000110100100000000000000000000000100001100000101100000",  -- ROS word 347
   "0000000101000010111110000000000000100000000000001000100100000011010011111100000000000001110100000000",  -- ROS word 3c4
   "0000001110100000011110000110011000000010000000000111100000000011110001001100000000000111010011100000",  -- ROS word 3c5
   "0000001101000010111110000000000000000000000000000000100010110100101101001111110100000110000011110000",  -- ROS word 3c6
   "0000000000000111011101000101101000000000000000000010100110000110101100010100000000000010000000000000",  -- ROS word 3c7
   "1000001101001100011110000001010000000001001000000100100010000011011011001100001100000111001111000000",  -- ROS word 444
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 445
   "1000000000000010111100000001010000000001001000001000100110000111011111001100000000000010000111000000",  -- ROS word 446
   "0000000000010010000000000110011000000011010000001101001010010100000000000000001000000000000000000000",  -- ROS word 447
   "1000000000000111111110000000000110010000000101010010100000000100011010000010110000000000110000110000",  -- ROS word 4c4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4c5
   "0000000000110111100010000101001000000011010000010010100000000000000010000000000000111100000000000000",  -- ROS word 4c6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 4c7
   "1000000000000111100010000000000000000000000000110010000100000110000100000000000000000000110000100000",  -- ROS word 544
   "1000000011000000000010000001111000000000000000001001011000000000000000000000000000000100000100000000",  -- ROS word 545
   "0000000000000000000010000000000000000000000000010010011000000000000010000000000000000000000100000000",  -- ROS word 546
   "0000000011000000000010000001111000000000000101101110001110010000000100000000000000000000000100000000",  -- ROS word 547
   "1000000000000000000000000100110010010000000000001011100010000100000010000000000000000000000100000000",  -- ROS word 5c4
   "1000000001000010111110000000000000000000000000001011100000010101101111100100100000000010100001110000",  -- ROS word 5c5
   "1000000001000010100000000000000000000000000000001000011110000000000011100000000000000110100001110000",  -- ROS word 5c6
   "1000001010001010000010000000000000000000000000110000011100000100000000000000000000010100010100000000",  -- ROS word 5c7
   "1000000000000000001010000000100000000000000000001001001000000000000000000000000000000000000001000000",  -- ROS word 644
   "0000000110000000000010000000000000000000000000001100100100000100000000000000000100001000000101100000",  -- ROS word 645
   "0000000110000000000010000000000000000000000000001100100110000100000000000000000100001100000011100000",  -- ROS word 646
   "0000000110100000000000000000011000000001100000001100100100000000000000000000000100001100000101100000",  -- ROS word 647
   "0000000000100000001000000000011000000001110000001010011100000100000010000000000000000000000011100000",  -- ROS word 6c4
   "0000001000000010000000000000011000000001101000000111011100000100000010000000000000000100000101100000",  -- ROS word 6c5
   "1000000110000000000010000000000000000000000000001101100100000000000000000000000000000000000011100000",  -- ROS word 6c6
   "0000000110000000000010000000000000000000000000000101100110000000000000000000000000000000000101100000",  -- ROS word 6c7
   "1000000000000010001010000000000000000000000000001110100110000000000010000000000000000000000001000000",  -- ROS word 744
   "0000000000000010001000000101101000000001101000001011100110000000000010000000000000000000000001000000",  -- ROS word 745
   "1000000000000010000000000000000000000001111000001110100010000000000010000000000000000100000011010000",  -- ROS word 746
   "0000000000000010000000000000000000000001111000001110100010000000000000000000000000000000000011010000",  -- ROS word 747
   "1000000000000010000000000000000000000001111000001011100110000000000010000000000000000001000110000000",  -- ROS word 7c4
   "0000000000000010000000000000000000000001111000001011100110000000000010000000000000000001000010010000",  -- ROS word 7c5
   "0000000100001100011110000000000000000000000000000110011010000101101111001100100000011010011101110000",  -- ROS word 7c6
   "0000000100001100011110000110101000000000000000010001011110000000000011001100100000011010011101110000",  -- ROS word 7c7
   "1000000000000111111011101000000011100000000000000011101000000100000000000000000010000000000000000000",  -- ROS word 844
   "1000001010000001100011010000111011100000000000000011101000000100000000000000000010000000000000000000",  -- ROS word 845
   "1000000000000000000001100101011011100000000000000011101000000100000000000000000000000000000100000000",  -- ROS word 846
   "1000000000000100100010000101110000000000000000110011011000000000000000000000000000000100000100000000",  -- ROS word 847
   "0000000000000000000000000000000010110000000000000111000100000000000000000000000000000100000100000000",  -- ROS word 8c4
   "1000000000000000001010000000000000010000000000001001001000000000000000010100100000000000000000000000",  -- ROS word 8c5
   "0000000000000000010010000000100000000000000000001000000100000100000000000000000000000000000100000000",  -- ROS word 8c6
   "0000000000000000000010000000000000000000000000000101101000000100000000000000000000000000000100000000",  -- ROS word 8c7
   "0000000000000000000010000000000000000000000000001100011010000000000000000000000000000000000100000000",  -- ROS word 944
   "0000000110000000000010000000011000000000000000001001001000000000000000000000000000000001011111010000",  -- ROS word 945
   "0000000000000010000010000110111000000011011000010110101000000000000010000000000000110100010000000000",  -- ROS word 946
   "1000000000000010000010000110111000000011011000010110101000000000000010000000000000100100010100000000",  -- ROS word 947
   "1000001101001100011110000001010000000001001000000100100010000011011011001100001100000111001111000000",  -- ROS word 9c4
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 9c5
   "1000000000000010111100000001010000000001001000010011011010000111011111001100001100000011001111000000",  -- ROS word 9c6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9c7
   "0000000000000000011110000110111000000000000000010101000000000100000011110100000000000000000100000000",  -- ROS word a44
   "1000000000000000000000000010000000000000000000010101001010000000000000000000000000000000000100000000",  -- ROS word a45
   "1000000000000111100010000001000110010000000101001100011010000100000000000000000000000100000100000000",  -- ROS word a46
   "0000000000000010000000000110010000000000001000010101000010000000000010000000000000000000000001000000",  -- ROS word a47
   "1000000000000000000010000000000000000000000000010101001100010100000000000000000000000000000011100000",  -- ROS word ac4
   "0000000000000000000010000000000000000000000001010101100010000100000000000000000000000000000100000000",  -- ROS word ac5
   "0011010000100000000000000000000000001000011001010101100010000000000000000000000000000100000100000000",  -- ROS word ac6
   "0000000000000010000000000000000000000001111000010101100110000100000000000000000000000000100000000000",  -- ROS word ac7
   "1000000000000000000000000000000011010000000010010110011111001110000100000000000000000000000100000000",  -- ROS word b44
   "1000000000000000000010000000000000000000000101010110100010010000000000000000000000000100000100000000",  -- ROS word b45
   "0000000000000000000000000000000011010000000010010110011110000000000000000000000000000100000100000000",  -- ROS word b46
   "1000000000010111100010000000000000001011110000010111100000000000000010000000000000000100110100110000",  -- ROS word b47
   "1000000001000000000000000000000000000000000001010111100010000000010100000000000000111001011100000000",  -- ROS word bc4
   "1010001011100111000000000101101000001000000000010111100010000100000001101100000000000010000111100000",  -- ROS word bc5
   "1000000001000000000000000001001000000000000000010100100010000110100010000000000000000100000011100000",  -- ROS word bc6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word bc7
   "0000000001010000000000000110110000000101001000011001011010000100000010000000000000000100100110011000",  -- ROS word c44
   "0000000001010000000010000110010000000101001000011001011100000000000000000000000000000100100010001000",  -- ROS word c45
   "0000000001000000000000000110110000000000000000011000000100000000000010000000000000111101011100000000",  -- ROS word c46
   "1000000000000010011001100000000000001101010000011000000100000100000010000011100001000000000100000000",  -- ROS word c47
   "0000000001010000000000000001111000000011010010111001100010000100011100000000000000111000000000000000",  -- ROS word cc4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word cc5
   "1000000000000000000010000010001000000000000000011001100000000000000000000000000000000100000100000000",  -- ROS word cc6
   "1000000000000000000010000110011000000000000000011001100100000010001010000000000000000101011100001000",  -- ROS word cc7
   "1000100000100000000010000110110000000100111000011010100000000000011000000000000000000101011111010000",  -- ROS word d44
   "1000000000010111100010000110011000000011010101011010010100000000000000000000000000000000010000000000",  -- ROS word d45
   "0000100000100000011110000000000000000110001000011010100000000100000001101110110000000011011111010000",  -- ROS word d46
   "0000000000000010000000000000000000001100000000011010100100000000011000000000000000000001011000000000",  -- ROS word d47
   "1000001011000111000010000000000000000000000000011011100010000110001001001111110000000010000001000000",  -- ROS word dc4
   "0000000001100111000000111000000000000100101000011011100000000000000000000011100001000000000011100000",  -- ROS word dc5
   "0000000000000111000000000000000000000000000000011011100010000100000010000011110000000100000100000000",  -- ROS word dc6
   "0000000001000000000000000000000000000000000000011011100000000000000010000000000000000101000111100000",  -- ROS word dc7
   "0000000000010010000000000000000000001100100000011100100100000000000000000000000000000000010000011000",  -- ROS word e44
   "0000000000000111100010000000000000000000000100111100100100000100000010000000000000000000110100110000",  -- ROS word e45
   "1000000000000010000000000001000000001100100000011100100000000100010100000000000000000000100111100000",  -- ROS word e46
   "1000001010000000000010000100111000000000000000111100000000000000010101001000100000000100000101000000",  -- ROS word e47
   "1010100000000110000010000110110000000000000000011101100101011000000000000000100001000000000001000000",  -- ROS word ec4
   "0010100000000110000010000110110000000000000100111101100101011000000010000000100001000100000001000000",  -- ROS word ec5
   "0011100000000111000010000000000000000000000011011101100010000100000011101100100001000110000000000000",  -- ROS word ec6
   "1000000000000010011000000110110000000000000000011101100110000100000000000000000000000101101000110000",  -- ROS word ec7
   "0000000000001011100010000000000000000000000000011110011010000000000000000000000000000000000100000000",  -- ROS word f44
   "0000000000000000000010000000000000000000000100111110100010000100000000000000000000000000000100000000",  -- ROS word f45
   "1000000000000000000010000000000000000000000001011110100100100000000000000000000000000100000100000000",  -- ROS word f46
   "1000000000000000011100000000000000000000000000011110100110000010001111000100000000000000000100000000",  -- ROS word f47
   "1000001001000010000001010000000000001110010000011111001010000010001000000000000000000000000100000000",  -- ROS word fc4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fc5
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fc6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fc7
   "1000001110000000011110000000000000000000000000000000100100111100101101001110110100000011110000000000",  -- ROS word 048
   "0000000100000000011110000000000000000000000000000000100100111100101101001110110100000011010100000000",  -- ROS word 049
   "1000000101000010111110000000000000100000000000010011100010000011010010000001100000000001110011000000",  -- ROS word 04a
   "1000000101000010111110000001001000100000000000001000100010000011010010000001100000000001110011000000",  -- ROS word 04b
   "1000000100000000000000000000000000000000000000000001100010000100000000000000000000000101110000000000",  -- ROS word 0c8
   "1000000001000010011100000001111000000000000000000001100000000011110111001110000000000110000000000000",  -- ROS word 0c9
   "0000000000000010111100000000000000000000000000000001100100000011011111001110111010000010000011110000",  -- ROS word 0ca
   "1000000000000000011100000010010000000000000000010011010010000000000000000000000000000000000100000000",  -- ROS word 0cb
   "1000000101000000000010110110011111100000000000000010100100000100000010000000000100000000101000000000",  -- ROS word 148
   "1000000101000000000010110000000111100000000000000010100110000000000010000000000100000000101000000000",  -- ROS word 149
   "1000000101010000000000110000000111100001010000000010100100000000000010000000000100000100101000000000",  -- ROS word 14a
   "1000000101000000000010110000000111100000000000000010100100000100100000000000000100000000101000000000",  -- ROS word 14b
   "1000000001000000000000000000000000000011011000000010100010000000101100000000000000000100000001000000",  -- ROS word 1c8
   "0000000000010000000001000110011000000001000000000011100010000011110110000000000000000100000100000000",  -- ROS word 1c9
   "1000000000000010111100000000000000000000000000000011100100000011011111001110111010000110000011110000",  -- ROS word 1ca
   "0000000000000010001010000000000000000001001000010011010010000100000010000000000000000000000100000000",  -- ROS word 1cb
   "1000000000000011000000000101000000000001011000010010010010000000111001001100000000000010000100110000",  -- ROS word 248
   "0000000000000010000000000000000000000001111000001000001000000000000010000000000000000001011000000000",  -- ROS word 249
   "0000000000000010111100000000000000000001001000000100100100000011011111001110111010000010000011110000",  -- ROS word 24a
   "0000000000000000011100000001000000000001011000010011100110100100000001001111110000000110000100000000",  -- ROS word 24b
   "0000000000000010001010000010110011100001111000000101100100000100000000000000000000000000101100000000",  -- ROS word 2c8
   "0000000000000010000000110010110011100001111000000101100100000100100000000000001010000100101100000000",  -- ROS word 2c9
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 2ca
   "0000000000000010000000110010110011100001111000000101100100000100100000000000001010001100000111100000",  -- ROS word 2cb
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 348
   "0000000000000010000000110000011000000001111000000110100100000000100000000000000100001000000011100000",  -- ROS word 349
   "0000000000000010001010110000011000000001111000000110100100000000000000000000000100001100000011100000",  -- ROS word 34a
   "0000000000000010000000110000000000000000000000000110100100000000000010000000000100001000000011100000",  -- ROS word 34b
   "0000000101000010111110000100100000100000000000001000100100000011010010000001100000000000000111110000",  -- ROS word 3c8
   "0000001110010010011100000110011000000011010000000111100000000011110001001100000000000111010100000000",  -- ROS word 3c9
   "1000001110000000011110000000000000000000000000000000100100111100101101001110110100000011110000000000",  -- ROS word 3ca
   "0000000101000010111110000000000000100000000000001000100010000011010011111100000000000001110111000000",  -- ROS word 3cb
   "1000000000000010111110000001011000000001001000000100100100000011011111001110111010000010000011110000",  -- ROS word 448
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 449
   "1000000000000000011100000000000000000001001000001000100110000111011111001100000000000010000100000000",  -- ROS word 44a
   "0000000000000010000000000000000000000000000000000110001110000000000000000000000000000001011000000000",  -- ROS word 44b
   "1000001010000000000010000000000000000000000100010010001000000000000010000000000000110000010000000000",  -- ROS word 4c8
   "1000000000000111000010101110010000000000000011001001100000001100000101011100000000000100000100000000",  -- ROS word 4c9
   "0000000000000000000010000001001000000000000101101100101000010000000010000000000000000000000100000000",  -- ROS word 4ca
   "0000000000000000000010000000000000000000000101101100101000010000000010000000000000000000000100000000",  -- ROS word 4cb
   "0000001010000000000010000000000000000000000100010001001100000000000010000000000000110100010000000000",  -- ROS word 548
   "1000000000000111000010100110000000000000000011001010100100000011000101100000100000000000000000000000",  -- ROS word 549
   "1000000011000000000000000000000101100000000101110000010110010000000010000000000000000000000100000000",  -- ROS word 54a
   "1000000000000000000000000000000101100000000101100000011000010000000010000000000000000000000100000000",  -- ROS word 54b
   "1000000000000010111100000000000000000000000000000111011110000000000010000000100000000100100001110000",  -- ROS word 5c8
   "1000000000000010111100000000000000000001111000001010001000000000000010000000100000000100100001110000",  -- ROS word 5c9
   "1000000000000000001000000010100000000000000000001011100110000000000010000000000000000000000100000000",  -- ROS word 5ca
   "1000000000000000001000000010100000000000000000001011100110000000000010000000000000000000000100000000",  -- ROS word 5cb
   "1000000000000010001010000000100000000001101000001101011100000100000010000000000100000100111101100000",  -- ROS word 648
   "0000000000000000000010000010010000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 649
   "1000000000000010000000000000011000000001111000000111011110000000000000000000000000000000101100000000",  -- ROS word 64a
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 64b
   "1000001000000010000000000000011000000001101000000000011100000100000010000000000000000000101100000000",  -- ROS word 6c8
   "0000000000000000000010000000000000000000000001001111011100000000000010000000000000000000000100000000",  -- ROS word 6c9
   "1000000110010000000010000000000011100001100000000101100110000100000010000000000000001000101001100000",  -- ROS word 6ca
   "1000000001000000000000000000000000000000000000001111011100000100000010000000000100000000111101100000",  -- ROS word 6cb
   "0000000000000111100010000000000000000000000000001110001000000010000100000000000000000100110000100000",  -- ROS word 748
   "0000000000000111100010000000000000000000000000001001100100000000000000000000000000000100000000100000",  -- ROS word 749
   "1000000000000111100000000001000000000000000000001110100100000000000010000000000000000100110000100000",  -- ROS word 74a
   "1000000111000000000010010000000000000000000000001100000110100000000000000000000000000001011000000000",  -- ROS word 74b
   "0000000000000000000000000110001000000000000000001000011110000100000000000000000000000100000100000000",  -- ROS word 7c8
   "0000001011000000000000000000000000000000000000001010010001001000000000000000000000000000000001000000",  -- ROS word 7c9
   "0000000000000111000010000000000000010001111000010000001110000000000011001100000000000010000100000000",  -- ROS word 7ca
   "1000000000000111000010000011010000000000000011001011100110000000000011001100000100000000010010100000",  -- ROS word 7cb
   "1000000111000000011110000000010101010000000000001010011110000100000011001100000000001111110100000000",  -- ROS word 848
   "0000000111000000011100000000000101010000000000001100000100000000000011001100000000001111110100000000",  -- ROS word 849
   "1000000110000000011110000000000101010000000000001100000010100000100101001100000000001111110100000000",  -- ROS word 84a
   "1000000111000000011100000000000101010000000000001100000100000000000001001100000000001011110100000000",  -- ROS word 84b
   "1000001101000000011000000000000000000000000000000100000010000100000011110100000100000110100000000000",  -- ROS word 8c8
   "1000001101000000011000000001001000000000000000000100000010000100000011110100000100000110100000000000",  -- ROS word 8c9
   "0000000000000111100010101000000000000011011000001100101010011000000010000000000000000100110000100000",  -- ROS word 8ca
   "0000000000000010000010001000000000000001111000001000000100000001000010000000000000000101011000000000",  -- ROS word 8cb
   "1000000110000000000000000000000011010000000000000110101000000100000010000000000000010100110000000000",  -- ROS word 948
   "1000000000000010000000000000011000110000000000001001001000000000000000000000000000000001011111010000",  -- ROS word 949
   "1000000000000010000000000000011000110001111000001001001000000000000000000000000000000001011111100000",  -- ROS word 94a
   "1000000000000010000000000000011000110001111000001001001000000000000000000000000000000001011111010000",  -- ROS word 94b
   "0000000000000011000000000101000000000001011000010011010010000000111001001100000000000110000100110000",  -- ROS word 9c8
   "1000000101000000011110010000000101000000000000000001100110000010000011001100000000000110101100000000",  -- ROS word 9c9
   "1000000000000111000000000101011000000000000000001111000110000100000010000000110000111100000000000000",  -- ROS word 9ca
   "1000000000000000000010000000000000000000000000010011010010000100000000000000000000000100000100000000",  -- ROS word 9cb
   "1000000000000000011100000011101000000000000000110100100100000010001001001111110000000010000100000000",  -- ROS word a48
   "0000000000000000000010000011110000000000000000010101000010000100000000000000000000000000000100000000",  -- ROS word a49
   "1011010000101000000010000100001000001000011000010101001000010100000000000000000000000100000100000000",  -- ROS word a4a
   "1000000000000010000010000000000000000000001000010101100000000100000000000000000000000000000001000000",  -- ROS word a4b
   "1000000000000000011100000000000000000000000001010101100110000000000100000000100000000100000000000000",  -- ROS word ac8
   "0000000000001111000010000000000000000000000000010101100100000100001100000000000000000100000011100000",  -- ROS word ac9
   "0000000000000000000010000000000000000000000000010101100110000100000000000000000000000000000100000000",  -- ROS word aca
   "1000000000000000000010000000011000000000000000000000011010000100000000000000000000000100000100000000",  -- ROS word acb
   "1000000000000101000010000000000000000000000001010110100100000100000010000000000000000100000100000000",  -- ROS word b48
   "0000000000000000000010000000000000000000000010110110011110000100000000000000000000000100000001000000",  -- ROS word b49
   "0000000000000111000000000000000000000000000011010110011110000100000001001100000000000110000100000000",  -- ROS word b4a
   "0000000000000000000010000000000000000011101000010110011110000100000000000000000000000100000011100000",  -- ROS word b4b
   "0000000001000000000000000111111000000000000000010111011110000101101000000000000000111101011100000000",  -- ROS word bc8
   "0000000000000000000000000100011000000000000000010111011110000100000010000000000000000100000100000000",  -- ROS word bc9
   "1000000001000000000000000111111000000000000000010111011110000101101000000000000000000100000011100000",  -- ROS word bca
   "1000000001000000000000000111111000000000000000010111011110000101101000000000000000000100000011100000",  -- ROS word bcb
   "1000000000000011000000000101101000001101000000011001000100000000000001110100000000000110000000110000",  -- ROS word c48
   "0000000000000011000001100101101000001101000000011001000100000000000000000011100001000100000100110000",  -- ROS word c49
   "1000000001000111000010000110011000000000000000011000100100000100000011001100000000000100000101000000",  -- ROS word c4a
   "0000000000000111100010100100101000000011011101011000100010000110100000010110100001000010110100110000",  -- ROS word c4b
   "0000000000000000000000000111011000000000000000011001100110000011111010000000000000000100000100000000",  -- ROS word cc8
   "0000000000000010000000000000000000000000000000011000010110000100000000000000000000000100000101001000",  -- ROS word cc9
   "0000001010000111100010000101101000000000000100011000101010000100000010000000000000110100010000000000",  -- ROS word cca
   "1000001010000111100010000101101000000000000100011000101010000100000010000000000000100100010100000000",  -- ROS word ccb
   "0000000001100000000010000110011000000110000000011010100010000100000000000000001110000101000011100000",  -- ROS word d48
   "0000001011100000000010000000000000000110000000011011001000000000000010000000000000000100000011100000",  -- ROS word d49
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d4a
   "1000000000010111100010000000000011010100001000011010100110000010000100000000000000000100000100000000",  -- ROS word d4b
   "0000000000000010000000000101111000001100010000011011100100000000000010000000000000000000010000000000",  -- ROS word dc8
   "0000001010000010000010000001111000001100111011011011100100000100000000000000000000000001101101000000",  -- ROS word dc9
   "1000000001000111000010000110110000000000000101011011100100000100000010000000000000011100000100000000",  -- ROS word dca
   "1000001011000111000010000110011000000000000011011011100110000000000000000000000000000000001000000000",  -- ROS word dcb
   "0000000000000111100000011001000000000000000111011100100110000010001010000000000000000100110100110000",  -- ROS word e48
   "0000000000000111100010000001001000000000000100111100100100000100000010000000000000000000110100110000",  -- ROS word e49
   "1000000000000010000000011110111000010000000000011100001100000100000000000010000000000100000000110000",  -- ROS word e4a
   "0000000000010010000000011000000000001100100000111100101000010110001010000000000000110000010000011000",  -- ROS word e4b
   "0000000000000000000010011000000000000000000101011101100010000100000000000000000000011000000100000011",  -- ROS word ec8
   "1000000000000000000010011000000000000000000000111101100110000000000000000000000000011100000100000011",  -- ROS word ec9
   "0000000000000000000010000000000000000000000101011101100010000100000000000000000000000000000100000000",  -- ROS word eca
   "1000000000000000000010000000000000000000000000111101100110000000000000000000000000000100000100000000",  -- ROS word ecb
   "1001010000001010000010000000000000000000000000011110100010000000000000000000000000000100000100000000",  -- ROS word f48
   "0010100000000000000010000000000000000000000000011110101000000110001000000000100001000000000100000000",  -- ROS word f49
   "0001010000001010000010000000000000000000000000011110101010000000000000000000000000000000000100000000",  -- ROS word f4a
   "0000000000000000000010000000000000001100101000011001101000010100000000000000000000000000000100000000",  -- ROS word f4b
   "1000000000000010000010000000000000001100100000011000010100000000000010000000000000000000010000000000",  -- ROS word fc8
   "0000000000000010000010000000000000001100100000011000010100000000000010000000000000000000010111100000",  -- ROS word fc9
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fca
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fcb
   "0000001110000000011110000000000000000000000000000000100110111100101101001110110100000111110000000000",  -- ROS word 04c
   "1000000100000000011110000000000000000000000000000000100110111100101101001110110100000111010100000000",  -- ROS word 04d
   "0000000101000010111110000000000000100000000000001000100000000011010010000001100000000101110011110000",  -- ROS word 04e
   "0000000101000010111110000001001000100000000000001000100000000011010010000001100000000101110011110000",  -- ROS word 04f
   "1000000101000000011110000001111101010000000000000001100110000101101111001100000000000111100100000000",  -- ROS word 0cc
   "1000000101000000011110000110101101010000000000010011100100000000000011001100000000000111100100000000",  -- ROS word 0cd
   "1000000101000111000010010110011101000011011000001111000000100000101101001100000000000110101100000000",  -- ROS word 0ce
   "1000000101000111000010010110110101000000000000010000011110000100000001001100000000000110101100000000",  -- ROS word 0cf
   "1000000101000111000000000001100000000000000000001101011110000100000000000001010100000100101000000000",  -- ROS word 14c
   "1000000101000000000010110000000111100000000000000010100110000001000000000000000100000000101000000000",  -- ROS word 14d
   "0000000101000000000000000110100101000000000000000100100110000000111000000000000000000000101001110000",  -- ROS word 14e
   "1000000101000111011110000000000000000000000000001111000100000000000001001111110100000011100011110000",  -- ROS word 14f
   "1000000101000000011100110000000111100000000000000010100100000000101101001110000000000110000000000000",  -- ROS word 1cc
   "1000000001010010000011000110011000000001010000000011100010000011110110000000000000000100000100000000",  -- ROS word 1cd
   "0000000000000010111100000000000000000000000000000011100110000011011111001110111010000010000011110000",  -- ROS word 1ce
   "0000000000000010001010000000000000000001001000010011010010000100000010000000000000000000000100000000",  -- ROS word 1cf
   "0000000101000000011100000001000101010000000000010011100100000000000010000000000000000101100100000000",  -- ROS word 24c
   "1000000101000000011100000010101101010000000000010011100101110000000010000000000000000001100100000000",  -- ROS word 24d
   "1000000000100000000000000000000010000011010000001111011110000100000000000000000000000000000100000000",  -- ROS word 24e
   "0000000000100000000000000000000010000011010000001110011110000100000000000000000000000100000100000000",  -- ROS word 24f
   "1000001000000010000000000000011000000001101000000111000010000100000000000000000000000000101100000000",  -- ROS word 2cc
   "0000001001000000000010000000000000000000000010001001000100000000000010000000000000000000000100000000",  -- ROS word 2cd
   "1000000000000000000010000000000000000000000000010001100010000110000110000000000000000100000100000000",  -- ROS word 2ce
   "1000000000000010000000000000100011100000000000000000101001001100000000000000000000000000101100000000",  -- ROS word 2cf
   "0000000000000010000000000000011000000001111000000110100100000000000000000000000000000100101100000000",  -- ROS word 34c
   "0000000000000010000000110000011000000001111000000110100100000000100000000000000100000000101000000000",  -- ROS word 34d
   "0000001011000000000000000000000000000000000000000110100110000100000010000000000000000000000001000000",  -- ROS word 34e
   "0000000001000000000010110110001000000000000000001001101001001100001110000000000000000100000011100000",  -- ROS word 34f
   "0000000101000010111110000100100000100000000000001000100100000011010010000001100000000000000111110000",  -- ROS word 3cc
   "0000000000000000001000000000000000000011101000000110010100000100000010000000000000000100000100000000",  -- ROS word 3cd
   "0000001110000000011110000000000000000000000000000000100110111100101101001110110100000111110000000000",  -- ROS word 3ce
   "1000000101000010111110000000000000100000000000001000100000000011010011111100000000000101110111110000",  -- ROS word 3cf
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 44c
   "1000000000000101000010000000000000000001111001001000001000000000000010000000000000000100000100000000",  -- ROS word 44d
   "1000000000000011000000000101000000000001011000010010010010010100111001001100000000000010000100110000",  -- ROS word 44e
   "1000000000000000001010000001000000100001011000010011100110100100000000000000000000000100000100000000",  -- ROS word 44f
   "0000000000000000000010000000000000000000000000001111001000010100000000000000000000000000000100000000",  -- ROS word 4cc
   "1000000011000000000000000111001011010000000000001101101000000000000000000000000000000000000100000000",  -- ROS word 4cd
   "0000000000000000000010000000000000000000000000010010011000000000000010000000000000000000000100000000",  -- ROS word 4ce
   "1000000011000000000000000111001011010000000101101100101000010000000010000000000000000000000100000000",  -- ROS word 4cf
   "1000000000000111100010000000000000000011011101001011000010000000000010000000000000000000000000100000",  -- ROS word 54c
   "1000000011000000000010000001111000000000000000001010011000000000000000000000000000000100000100000000",  -- ROS word 54d
   "1000000000000111100010000000000000000000000101001011000010000000000010000000000000000000000000100000",  -- ROS word 54e
   "0000000011000000000000000001111101100000000101101100010110010000000010000000000000000100000100000000",  -- ROS word 54f
   "0000000000000000000010000010010000000000000000001011100110000000000010000000000000000000000100000000",  -- ROS word 5cc
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 5cd
   "1000001011000000000000000000000000000000000000001011100110000100000010000000000000000100000001000000",  -- ROS word 5ce
   "1000000001000000000010100110000000000000000011001001100100000011000100011110110000000000000011100000",  -- ROS word 5cf
   "0000000000001010000010000000000000000000000110101101011000000100000000000000000000000000000100000000",  -- ROS word 64c
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 64d
   "0000000000000010000000000000011000000001111000000000011110000000000000000000000000000100101100000000",  -- ROS word 64e
   "0000000000000000000010000000000000000000000000000010101000000000000000000000000000000000000100000000",  -- ROS word 64f
   "1000000000000111000000000110110000000000000011001101100110000000000011001100000000000010000100000000",  -- ROS word 6cc
   "1000000000000111111100000001111000000000000000001110101010000000000001101000000000011100000000110000",  -- ROS word 6cd
   "0000000110100000000010000000000000000001110000001001011100000100000010000000001010000001001100000000",  -- ROS word 6ce
   "0000000000000111100010000000000000000000000000101110101010000000000000000000000000000000110100110000",  -- ROS word 6cf
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 74c
   "1000000000000010000010000101101000000001101000001011100110000000000010000000000000000000000011010000",  -- ROS word 74d
   "0000000000000000000010000011110000000000000000000000001000000000000000000000000000000000000100000000",  -- ROS word 74e
   "1000000000001011000000000000000000000000000001001110100110000100000001001100000000000100000000000000",  -- ROS word 74f
   "1000000101000000011110000000000011010000000000001001100010000000000001110011101010000101100111110000",  -- ROS word 7cc
   "1000000101000000011110000000000011010000000000001111100110000100011011111001110000000001100001010000",  -- ROS word 7cd
   "0000000000010000000010111000000000000010111000001111100110000100000000000000000000000100000001000000",  -- ROS word 7ce
   "0000000101000000011100111000000000000010011000001111100110000100000011100000100100000000101001110000",  -- ROS word 7cf
   "0000000000000010000000000000000000000000000000001101011110000100000010000000000000000000000001000000",  -- ROS word 84c
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 84d
   "1000000000000000001000000010010000000000000000001011100110000000000010000000000000000000000100000000",  -- ROS word 84e
   "1000000000000000001010000000000000000001101000001001011110000100000010000000000000000100000100000000",  -- ROS word 84f
   "0000001001000101000000001000000000000001111101010001100100000100000010000000000000000100000100000000",  -- ROS word 8cc
   "1000001001000101001010001000000000000001111000000100100100000000000010000000000000000100000100000000",  -- ROS word 8cd
   "0000000000000100011100001000000000000001111101001001010100000100000010110100000000000110000100000000",  -- ROS word 8ce
   "0000000000000100000010001000000000000001111101001000100110000000000010000000000000000000000100000000",  -- ROS word 8cf
   "0000001001000000000000000001000000000000000000010000001010000000000000000000000000000001000000000000",  -- ROS word 94c
   "1000001001000000000010000001001000000000000000010000001010000000000000000000000000000001000000000000",  -- ROS word 94d
   "1000000110000010000000000000011000000001111000001001001000000000000000000000000000000001011111100000",  -- ROS word 94e
   "1000000110000010000000000000011000000001111000001001001000000000000000000000000000000001011111010000",  -- ROS word 94f
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 9cc
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9cd
   "0000000000000011000000000010010000000001011000010011100110000000000001001100000000000110000100000000",  -- ROS word 9ce
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 9cf
   "1000000000000000000000000110001000000000000001010100100110000000001110000000000000000000000100000000",  -- ROS word a4c
   "0000000000010010000000000011110000000001110000010101000100000100110110000000000000000001011000000000",  -- ROS word a4d
   "1000000000000000000010000000000000000000000000010100101000000010000010000000000000000100000100000000",  -- ROS word a4e
   "1000000000000000000010000000011000000000000000010100101000000010000010000000000000000100000100000000",  -- ROS word a4f
   "1000000000000111000000000000000000000000000000110101100100000010001011001111110000000010000100000000",  -- ROS word acc
   "0000000000000000011110111000000000000000000000010101100111000000000000000000000000000000000100000000",  -- ROS word acd
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word ace
   "1000000000000000000010000000000000000000000001010101010110000100000000000000000000000100000100000000",  -- ROS word acf
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word b4c
   "0000000000000000000010000000011000000000000000010101100100000000000000000000000000011000000100000000",  -- ROS word b4d
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word b4e
   "1000000000000010011100000000000000000000001001010111000010000000000010000011110000000000000100000000",  -- ROS word b4f
   "1000000000000010000000000000000000000000000000010111100110000100000000000000000000000100000001000000",  -- ROS word bcc
   "0000000000000010000000000000000000000000000000010111100110000100000010000000000000000000000001000000",  -- ROS word bcd
   "1000000000000000000010011000000000000001111000010111101010000000000000000000000000000001000000000000",  -- ROS word bce
   "0000000000000000000010000000000000000001111000010111101000000000000010000000000000000000000100000000",  -- ROS word bcf
   "0000000000000101000001000000000000000011011000011000100110000100000001001010100001000110000100000000",  -- ROS word c4c
   "1000000000100111111100000111011000000101000000011000100110000100000010000000100000000000000100001000",  -- ROS word c4d
   "1000000000010010000011000110001000000101011000011000100001011110001000000000000000000001000000000000",  -- ROS word c4e
   "1000000000000111000010000000000000001101000000011000101010000100000000000000110000000100000100000000",  -- ROS word c4f
   "1000000000100000000000000000000000100101001000011011000000000100000010000000000000010100000000000000",  -- ROS word ccc
   "0000000000100000000000000000000000100101001000011011000000000100000000000000000000010000000000000000",  -- ROS word ccd
   "1000000000000000000000000000000000100000000000011011000110000100000010000000000000010100000000000000",  -- ROS word cce
   "0100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word ccf
   "0000000000000000000010000111011000001100001000011010100110000100000000000000000000000000000100000000",  -- ROS word d4c
   "0000000001100000000000000110010000000100001000011010101000000000000000000000000000000000000011100000",  -- ROS word d4d
   "1000000000000010000000000110010000001100010000011010011000000000000010000000000000000101000000000000",  -- ROS word d4e
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d4f
   "0000000000000011100010000110100000001100011000011011100110000000000010000000000000000101101000110000",  -- ROS word dcc
   "0000000000010000000000000110100000000100101000011011100110000101011010000000000000000100000100000000",  -- ROS word dcd
   "0000001010010000011011001110100000000100100000011011101000000110001010000011100001000100000001000000",  -- ROS word dce
   "0000000000100000000000000110011000000101011101011011010000000100000010000000000000111000000000000000",  -- ROS word dcf
   "0000000000010000000010000000000000000100110010011100001010000100000000000000000000000000000100000000",  -- ROS word e4c
   "1000001011001111010100110000000000000000000000011101001111010100000000000010100001110100000000000000",  -- ROS word e4d
   "0000000000000000000010000001001000000000000000011100011110000011111010000000000000000000000100000000",  -- ROS word e4e
   "1000000000000010000010000000000000001100100000011100011100000100010100000000000000000000010000000000",  -- ROS word e4f
   "0011100000000111000010000000000000000000000101011101100110000000000011101100100001000110000000000000",  -- ROS word ecc
   "1001010000001010000010000000000000000000000011011101100010000100000010000000000000000100000100000000",  -- ROS word ecd
   "1000000000011111000000000000000000000100111000011101011000000001011010000000000000000100000000001011",  -- ROS word ece
   "1000000000000111110100100110101000001100011000011101100000000000001111010000100001000100000001000000",  -- ROS word ecf
   "1010100000000111100000000101011000001100100000011110000010000010001010000000100001000100000001000000",  -- ROS word f4c
   "0000000000000000011010000000000000000000000000011110100110000000000000000011110000000000000100000000",  -- ROS word f4d
   "1000000000000010000000000000000000000000000000011110100110000100000010000000000000000001101101000000",  -- ROS word f4e
   "1000000000100111100010000000000000000101001101011011001100000000000000000000000000000100010111100000",  -- ROS word f4f
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fcc
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word fcd
   "1000000000110000000000011000000000000110111000011111010110000000000000000000000000111100000000000000",  -- ROS word fce
   "1000000000110000000000011000011000000011010000011111010110000000000000000000000000111100000000000000",  -- ROS word fcf
   "1000001100000000000010000000000000000000000000000000101000000000000010000000001010000000000001000000",  -- ROS word 050
   "0000000000000010000000110010110011100001111000000000101010000000100000000000001010001101001111100000",  -- ROS word 051
   "1000000000000000001000000101000000000001111000001001001000000000000000000000000000000000000100000000",  -- ROS word 052
   "1000001001000000000010000000000000000000000001010001001010000000000000000000001000000000000000000000",  -- ROS word 053
   "1000000000000101100010000100110000000000000000001101011000000000000010000000000000000100000100000000",  -- ROS word 0d0
   "1000000001100000000010000111011101100010010100000001101000000100000000000000000000000000000011100000",  -- ROS word 0d1
   "1000000000000011000010000000000000000000000000001110011000000010000100000000100000000000000000110000",  -- ROS word 0d2
   "1000000000000000011100000000000000000000000000100111000000000000011110000010110000000100000000000000",  -- ROS word 0d3
   "1000000000000100100000000000000011010000000000000000001001100000000000000000000000000000000100000000",  -- ROS word 150
   "1000000000000100100010000000000000000000000110100011101000000000000010000000000000000100000100000000",  -- ROS word 151
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 152
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 153
   "0000000000000100100010000000000000000000000110101101011000000100000000000000000000000000000100000000",  -- ROS word 1d0
   "1000000000001111011000000000000011100000000000001101011000000100000000000000000010000100000000000000",  -- ROS word 1d1
   "0000000000000000001000000000000000000000000000000011101000000000000000000000000000000100000100000000",  -- ROS word 1d2
   "1000000000001110101110000000000000000000000000001100000000000000000000000000000000000100000100000000",  -- ROS word 1d3
   "1000000000000000010000000000000000000000000000010000001110000100010100000000000000000000000100000000",  -- ROS word 250
   "1000000000000000000010000000000000000000000000000110010000000011011100000000000000000100000100000000",  -- ROS word 251
   "1000000000100000000111010111111000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 252
   "1000000000000010001010000000000000100001011000010011100110100100000000000000000000000100000100000000",  -- ROS word 253
   "1000000000000000000010000000000010100000000000000110011110000100000010000000000000000100000100000000",  -- ROS word 2d0
   "0000000000000000010000000000101010010000000000010000001110000100000010000000000000000100000100000000",  -- ROS word 2d1
   "1000000000000000000010000000000000000000000000000110011110000100000010000000000000000100000100000000",  -- ROS word 2d2
   "0000000000000000000010000000000010010000000110110001011000000100000010000000000000000000000100000000",  -- ROS word 2d3
   "0000000000000010000000000110111110010011011101110110101000000001010100000000000000110000010000000000",  -- ROS word 350
   "1000000000000010000000000110111110010011011101110110101000000001010100000000000000100000010100000000",  -- ROS word 351
   "1000000000000000000000000101001000000000000001001111000000000100000010000000000000000000000100000000",  -- ROS word 352
   "0000000000000111100010000100110110010000000101010010100010000000000000000000000000000100001000110000",  -- ROS word 353
   "1000000000000111100010000110011101110000000101000100000010000000000000000000000000100100010100000000",  -- ROS word 3d0
   "0000000000000111100010000110011101110000000101000100000010000000000000000000000000110100010000000000",  -- ROS word 3d1
   "0000000000000111100010000110011101110000000101000100000010000000000000000000000000110100010000000000",  -- ROS word 3d2
   "0000000000000111100010000110011101110000000101000100000010000000000000000000000000110100010000000000",  -- ROS word 3d3
   "1000000000000111000010110110001000000000000000001010101001001100001111110100000000000100000100000000",  -- ROS word 450
   "0000000000000111000000000000000000000000000000000110100110000110001111110100000000000100000100000000",  -- ROS word 451
   "1000000000000000000010000000000000000000000101101010100010010000000000000000000000000100000100000000",  -- ROS word 452
   "1000001011000000000000000000000000000000000101101010100010010000000000000000000000000100000001000000",  -- ROS word 453
   "1000000000000111000010101110010000000000000011001000101000001100000010111100110000000100000100000000",  -- ROS word 4d0
   "0000001010000000000010000000000000000000000100010010001000000000000000000000000000110100010000000000",  -- ROS word 4d1
   "1000000000000000000010101110010011010000000011001011000000001100000010000000000000000100000100000000",  -- ROS word 4d2
   "1000000000000000000010101110010011010000000011001011000000001100000010000000000000000100000100000000",  -- ROS word 4d3
   "0000000000000111000010101110010000000000000011001000101000001100000000111100110000000000000100000000",  -- ROS word 550
   "0000001010000000000010000000000000000000000100010010001000000000000000000000000000110100010000000000",  -- ROS word 551
   "1000000000000000000010101110010011010000000011001011000000001100000010000000000000000100000100000000",  -- ROS word 552
   "1000000000000000000010101110010011010000000011001011000000001100000010000000000000000100000100000000",  -- ROS word 553
   "0000000000000000000010000000000000000000000000001001100100000000000010000000000000000000000100000000",  -- ROS word 5d0
   "1000000000000100100010000000000000000000000000101001100100000000000010011110110000000100000100000000",  -- ROS word 5d1
   "0000000000000000000010000000000000000000000000001001100000000000000000000000000000000000000100000000",  -- ROS word 5d2
   "0000000000000100100010000000000000000000000000101001100000000000000010000000000000000000000100000000",  -- ROS word 5d3
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 650
   "0000000000000000000010000000000000000000000000001110100100010100000000000000000000000000000100000000",  -- ROS word 651
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 652
   "0000000000000000000010000000000000000000000000010010011000000000000010000000000000000000000100000000",  -- ROS word 653
   "0000000000000111000010101110010000000000000011001101101000001100000001011100000000000000000100000000",  -- ROS word 6d0
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 6d1
   "0000000000000000000010000000000000000000000101101100101000010000000010000000000000000000000100000000",  -- ROS word 6d2
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word 6d3
   "1000000000000111000000000000000000000000000000001010010110000010001110111100110000000000000100000000",  -- ROS word 750
   "1000001010000000000000000001001010000000000100010010001000000000000000000000000000110100010000000000",  -- ROS word 751
   "1000000000000000000010101110010011010000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 752
   "1000000000000000000010101110010011010000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 753
   "1000000000000111000010100110000000000000000011001010000100000011000100111100110000000100000100000000",  -- ROS word 7d0
   "1000001010000000000000000001001010000000000100010010001000000000000000000000000000110100010000000000",  -- ROS word 7d1
   "1000000000000000000010101110010011010000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 7d2
   "1000000000000000000010101110010011010000000011001111001000001100000010000000000000000100000100000000",  -- ROS word 7d3
   "1000001001000000000010000000000000000000000000001000011000000000000010000000000000000100000100000000",  -- ROS word 850
   "0000000001000000000000000000000000000000000000000110011000000000000010000000000000000000000011100000",  -- ROS word 851
   "0000001001000000000010000101101000000000000000010000001000100000000000000000000000000000000100000000",  -- ROS word 852
   "1000000000000000000010000000000000000000000101110010001000000100000010000000000000000100000100000000",  -- ROS word 853
   "1000001011000000000000000000000000000000000000010011000100000000010010000000000000000100000001000000",  -- ROS word 8d0
   "0000000000000000000010000000000000000000000000010011000100000100010010000000000000000000000100000000",  -- ROS word 8d1
   "1000001011000000000010000001000000000000000000010000101000010100010010000000000000000000000001000000",  -- ROS word 8d2
   "1000000000000000000000000001000000000000000000010000101000010100000000000000000000000000000100000000",  -- ROS word 8d3
   "0000000000000111100010000000000000000000000000001010000110000000000000000000000000000100110000100000",  -- ROS word 950
   "0000000000000000000010000000000000000000000000010010101000010000000000000000000000000000000100000000",  -- ROS word 951
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 952
   "1000000000000111000000101110000000000000000000010011001000001110001001001100000000000100000000000000",  -- ROS word 953
   "0000000000000011000000000101000000000001011000010011010010000000111001111100000000000110000100110000",  -- ROS word 9d0
   "1000000000100000000010000000000000000011010000010010001010101100000010000000000000000100000100000000",  -- ROS word 9d1
   "0000001101000010111110000000000000000000000000010011101010000000000001001110111010000111001011110000",  -- ROS word 9d2
   "0000000000000000001010000000000000000001011000010011010010000000000000000000000000000000000100000000",  -- ROS word 9d3
   "1000000000000000000000000011010000000000000000010101011000000101101110000000000000000000000100000000",  -- ROS word a50
   "0000000000000000000000000011010000000000000000010100101000000101101110000000000000000100000100000000",  -- ROS word a51
   "1000000000000010000000000000000000000000000000010100101010000101001110000000000000000100000001000000",  -- ROS word a52
   "0000000000000000000010000000000000000000000000010100101010000001001110000000000000000000000100000000",  -- ROS word a53
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word ad0
   "1000010000010000000010000101001000000011010000001111011010000100000000000000000000000100000100000000",  -- ROS word ad1
   "1000000000000000000000000101001000000000000000001101011000000100000010000000000000000000000100000000",  -- ROS word ad2
   "0000000000000000000000000100000000000000000000010110011000000100000000000000000000000100000100000000",  -- ROS word ad3
   "1000000110000000100000000101101101110000000010000110101000000110000100000000000000010100110000000000",  -- ROS word b50
   "1000000000110000000000000001111011011000010000110111010000000100000000000000000000000000000100000000",  -- ROS word b51
   "1000000000000001000000000000000000000000000000010110101010011100010100000000000000000000000100000000",  -- ROS word b52
   "0000000001100000000000000011001010110011010000010111000000101101010100000000000000011100000100000000",  -- ROS word b53
   "0000000000000100100010000000000000000000000001010110000100000000000000000000000000000000000100000000",  -- ROS word bd0
   "1000000000000000000010000000000000000000000000010111101010000101010000000000000000000100000100000000",  -- ROS word bd1
   "0000000000000000000000000101001000000000000000010111101000000100000010000000000000000100000100000000",  -- ROS word bd2
   "0000000000000000000010000000000010010000000000001101011000000100000010000000000000000000000100000000",  -- ROS word bd3
   "0000000000000111000000000110111000000010011011111000101000000000000011001100000000000100100100110000",  -- ROS word c50
   "0000000000111111000010000000101000000101101101011000011100000101011010000000000000000100000001000000",  -- ROS word c51
   "0000000000000110000010000100111000001101001101011000100100000010100011101100000000000010000101000000",  -- ROS word c52
   "1000000000000010011110000110110000001101010000011000101010000010100010110100000000000111011101000000",  -- ROS word c53
   "0000000000000000011011001000000000000000000000011101010110000000000000000011100001000000000100000000",  -- ROS word cd0
   "0000000000000111000010000000000000001101000000011001011111010100000010110100000000000010000100000000",  -- ROS word cd1
   "0000000001100000000000000000000000000100110000011000010110000100000010000000000000000001101001001000",  -- ROS word cd2
   "0000000000000111000010000101101000001101000000011001011110000100000010110100000000000010000100000000",  -- ROS word cd3
   "0000000001100000000010000110101000000100010000011010101000000000000010000000000000000101011011000000",  -- ROS word d50
   "0000001011010000000010000110101000000100100000011010101000000110101100000000000000000101000011000000",  -- ROS word d51
   "0000000000100000011100100000000000000101000000011010101010000110101100000000100001000000000001000000",  -- ROS word d52
   "1000000000100000011110000000000000000101000000011010101010000110101100000000000000000000000001000000",  -- ROS word d53
   "1000000000100000000000000110110000000100001000011011101000000000000010000000000000000000000100000000",  -- ROS word dd0
   "0000000000000111000011000110010000001110110000011011101000000100000000000000100001000000000100000000",  -- ROS word dd1
   "0000001011100111111100000001000000000100000000011011000010000100000001001000100000110100010100000000",  -- ROS word dd2
   "1000000000000000010100001110011000000000000000011101010100000100000010000010100001000100000000000000",  -- ROS word dd3
   "0000000000000010000010010000000000001100101111011100101010000100000010000000000000000000000100110000",  -- ROS word e50
   "0000001011001111010110010000000000000000000000011101001111010100000000000010100001110100000000000000",  -- ROS word e51
   "1000000000000010000000000000000000001100101111011100101010000100000010000000000000000000000100110000",  -- ROS word e52
   "1000001011001111010100100001000000000000000000011101001111010100000000000010100001110100000000000000",  -- ROS word e53
   "1000001001001011100010000000000000000000000000011101100000000000000001000100000000000010000000000000",  -- ROS word ed0
   "0000001001000000000010000000000000000000000000011101101000000100000000000000000000000000000100000000",  -- ROS word ed1
   "0001010000001010000010000000000000000000000001011101101000000100000010000000000000000000000100000000",  -- ROS word ed2
   "1000000000001011100010000000000000000000000000011101100000000000000001000100000000000010000000000000",  -- ROS word ed3
   "0000000001100000000000000110001000000100100000011111000010000000000010000000000000000000000000001000",  -- ROS word f50
   "0000000000000000000010000001001000000000000000011110011010000010001000000000000000000000000100000000",  -- ROS word f51
   "1000001010000000000000000010111010000000000000011110101010000000011010000000000000000100010001001000",  -- ROS word f52
   "0000000000000000000011010000000000000000000000011110100000010110001000000000000000000000000100000000",  -- ROS word f53
   "1000000000000000000000000110100000000000000000010110010110000000000010000000000000000000000100000000",  -- ROS word fd0
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word fd1
   "1000010000000000000000011000000000000000000000010110011110000000000000000000000000110000000100000000",  -- ROS word fd2
   "0000000000000111100010000000000000000000000101010110100100000000000000000000000000000000110100110000",  -- ROS word fd3
   "1000000000000010001010000000100000000001101000001001001000000000000000000000000000000001011000000000",  -- ROS word 054
   "1000001100000000000010000000000000000000000000000000101000000000000010000000001010000001011000000000",  -- ROS word 055
   "0000001101000111000010000000000000000000000000001001001000000110100011101100001000000010000100000000",  -- ROS word 056
   "1000001101000000000000000000000000000000000000010000011010000100000010000000001000000100000000000000",  -- ROS word 057
   "1000001001000010000000111110100000000000000000001011000100000111010000000000000000000101011000000000",  -- ROS word 0d4
   "0000001001000010000010111110110000000000000000001011000100000111010000000000000000000101011000000000",  -- ROS word 0d5
   "0000001010000000000010000101101000000000000000000001001000000000000000000000000000000100000001000000",  -- ROS word 0d6
   "1000000000010000000010000000000000000011010000001010001000000100000010000000000000000000000001000000",  -- ROS word 0d7
   "0000000000000111000000000110000000000000000000000010101010000000001111100000100000000000000000000000",  -- ROS word 154
   "0000000000000000000010000000000000000000000101000010101010000100000000000000000000000000000100000000",  -- ROS word 155
   "0000000000000000000000000101111000000000000000001001101010000000000010000000000000000100000100000000",  -- ROS word 156
   "0000000001000100100000000000000000000000000000010011001000000000000010000000000000000000000011100000",  -- ROS word 157
   "1000001101000000000000000000000000000000000000001010101010000000000000000000000000000000000100000000",  -- ROS word 1d4
   "1000000000000000000000000001001011010000000000001011101010000100000000000000000000000000000100000000",  -- ROS word 1d5
   "0000000000000000000000000001000001010000000000001011101010000000000000000000000000000100000100000000",  -- ROS word 1d6
   "0000001101000000000000000001001000000000000000001010101010000000000000000000000100011000110000000000",  -- ROS word 1d7
   "0000000000000000011100000000000000000011011000000100101010100000000010110100000000000110000100000000",  -- ROS word 254
   "1000000000010010000000000000000000000011010000000011101010000011001000000000000100000100111001000000",  -- ROS word 255
   "0000000000000000011100000000000000000011011000000100101010100000000010110111110000000110000100000000",  -- ROS word 256
   "1000000000000010000000000000000000000000000000000011101010000011001000000000000000000100000001000000",  -- ROS word 257
   "0000001101010010011100000000000000000011010000000100101010010100000001000100110100000110111101000000",  -- ROS word 2d4
   "0000001101010010011100000000000000000011010000000100101010010100000001000100110100000110111101000000",  -- ROS word 2d5
   "1000000000000111000000000110000000000000000000000110101010000000001111100000100000000100000000000000",  -- ROS word 2d6
   "1000000000000111000000000110000000000000000000000110101010000100001111110000100000000000000100000000",  -- ROS word 2d7
   "0000001101000111000010000110000000000000000000000110101010000000001111100000100000000100000000000000",  -- ROS word 354
   "1000000000000000011000000111000001010011011000000101101011011000000001001110110000000110000000000000",  -- ROS word 355
   "1000001101000111000010000110000000000000000000000110101010000100001111110000100100011000110000000000",  -- ROS word 356
   "1000000000000000011010000111000011010011011000000101101011011100000011001111110000000110000100000000",  -- ROS word 357
   "1000001101000000000000000000000000000011011000000101101010000000000000000000000000000000000100000000",  -- ROS word 3d4
   "0000000000000000000000000001001011010000000000000110101010000100000000000000000000000100000100000000",  -- ROS word 3d5
   "1000000000000000000000000001000001010000000000000110101010000000000000000000000000000000000100000000",  -- ROS word 3d6
   "0000001101000000000000000001001000000011011000000101101010000000000000000000000100011000110000000000",  -- ROS word 3d7
   "1000000000000101000000000111011000000000000000001000101010010100000010000000000000000000000100000000",  -- ROS word 454
   "1000000000000000011100000000000000000000000000001011000010000100000010000000100000000100000000000000",  -- ROS word 455
   "1000000000000100000000000000000000000000000000001000101010010100000010000000000000000000000100000000",  -- ROS word 456
   "1000000000000000011100000000000000000000000000001011000010000100000011001100100000000110000000000000",  -- ROS word 457
   "1000000000000000000010000000000000000011011000001000101010011000000000000000000000000100000100000000",  -- ROS word 4d4
   "1000001011000000000000000111001000000000000000000010101010000100000010000000000000000100000001000000",  -- ROS word 4d5
   "1000000000000000000010000000000000000011011000001000101010011000000000000000000000000100000100000000",  -- ROS word 4d6
   "0000000000000000000000000111000001010000000000000010101010000000000000000000000000000100000100000000",  -- ROS word 4d7
   "0000001101000000011100101101111000000011011101101010001010101100000001000100110100000110111101000000",  -- ROS word 554
   "0000001101000000011100101101111000000011011101101010001010101100000001000100110100000110111101000000",  -- ROS word 555
   "0000000000000111000000000110000000000000000000001011101010000000001111100000100000000000000000000000",  -- ROS word 556
   "0000000000000111000000000110000000000000000000001011101010000100001111110000100000000100000100000000",  -- ROS word 557
   "1000001101000111000010000110000000000000000000001011101010000000001111100000100000000000000000000000",  -- ROS word 5d4
   "1000000000000000011000000111000001010000000000001010101011011000000001001110110000000110000000000000",  -- ROS word 5d5
   "0000001101000111000010000110000000000000000000001011101010000100001111110000100100011100110000000000",  -- ROS word 5d6
   "1000000000000000011010000111000011010000000000001010101011011100000011001111110000000110000100000000",  -- ROS word 5d7
   "0000000000010010000000000000000000000011010000010001100100000100000000000000001010000000000001000000",  -- ROS word 654
   "0000000000000101000010000111011010000000000000001111000110000000000010000000000100000000000100000010",  -- ROS word 655
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 656
   "0000000000000100000010000000000010000000000000001111000110000000000010000000000100000000000100000010",  -- ROS word 657
   "0000000000000000011000000101111000000000000101101111010110000010001111001110111000000110000100000000",  -- ROS word 6d4
   "0000000000000111000000000110000000000011011000001110001010101100001111110000101010000000000001000000",  -- ROS word 6d5
   "1000000000010010011110000110011000000011010000001110010110000010001110110110111000000110000100000000",  -- ROS word 6d6
   "0000000000000111000000000110000000000011011000001110001010101100001111110000101010000000000001000000",  -- ROS word 6d7
   "1000000000000111000010110110100000000000000011001110101011001100101111001100000000000000000000000000",  -- ROS word 754
   "0000000000000000000010000000000000000000000101101101100110000100000010000000000000000000000100000000",  -- ROS word 755
   "0000000000000000000000000110010000000000000101110000010110101100000000000000000000000100000100000000",  -- ROS word 756
   "0000000000000000000000000110010000000000000101110000010110101100000000000000000000000100000100000000",  -- ROS word 757
   "0000000000000000000000011000000011010000000000001001010100000100000000000000001010000001001000000001",  -- ROS word 7d4
   "0000001101000000011110000000000000000000000000001111101010000100000010110100000100000010100100000000",  -- ROS word 7d5
   "1000000001000000000000000101101000000000000000001100000110000100000010000000000000000100000011100000",  -- ROS word 7d6
   "0000000000000000000010011000000000000000000000001111101010100000000000000000000000000100100000000000",  -- ROS word 7d7
   "1000001101000010011100000000000000000000000000001010101010000000000000110100000000000010000100000000",  -- ROS word 854
   "1000000000000010011100000001001011010000000000001011101010000100000000110100000000000010000100000000",  -- ROS word 855
   "1000000000000010011110000000000000000000000000001011101010000000000000110100000000000110000100000000",  -- ROS word 856
   "0000000000000000000010000010100000000000000000010010000110000100000000000000000000000000000100000000",  -- ROS word 857
   "0000000000000111100010000000000000000000000000010011000000000000000010000000000000000100000000100000",  -- ROS word 8d4
   "1000000000000111100010000000000000000000000000010011000000000000000000000000000000000000000000100000",  -- ROS word 8d5
   "0000000000000111100010000000000000000000000000010010001010000000000000000000000000000100000000100000",  -- ROS word 8d6
   "0000000000000111100010000000000000000000000000010010001010000000000000000000000000000100000000100000",  -- ROS word 8d7
   "0000000000000000000010000000000000000000000011010010101010000100000010000000000000000000000100000000",  -- ROS word 954
   "0000000000000000000010011000000000000000000000010011001100000100000000000000000000000100100000000000",  -- ROS word 955
   "1000000000000000011010000000000000000000000000010010101010101100000011110100000000000010000000000000",  -- ROS word 956
   "0000000000100000000010000000000000000011010000001110001100101101100100000000000000000000000100000000",  -- ROS word 957
   "1000000000000000000010000000000000000001001000010011101000000011011011001100000000000110000100000000",  -- ROS word 9d4
   "1000000101000000011100000000110000000000000000010010011110000100000000000001100100000000000101110000",  -- ROS word 9d5
   "1000000000100000000111010000000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word 9d6
   "0000001010001010000010000000000000000000000000010011101010000100000000000000000000010000010100000000",  -- ROS word 9d7
   "0000001010000000000000000010000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word a54
   "0000000000000000000010000000000000000000000000010101011000000000101110000000000000000000000100000000",  -- ROS word a55
   "0000001010000000000000000010000000000000000000010101001010000000000000000000000000000000000000001000",  -- ROS word a56
   "1000000000000000000000111000000000000000000101010110010000000010100010000000000000000000000100110000",  -- ROS word a57
   "1000000000000000011100000000000000000000000000010101101010110100110111001111110000000010000100000000",  -- ROS word ad4
   "0011000000100000000010000000000000001000000000010101100000000000000010000000000000000000000100000000",  -- ROS word ad5
   "1000000000001000000000000000000000000000000000010101001010010100000000000000000000000000000100000000",  -- ROS word ad6
   "0011000000100000000010000000000000001000000000010101100000000000000010000000000000000000000100000000",  -- ROS word ad7
   "1000000001000000000000000110011000000000000000010110101000000101101000000000000000111001011100000000",  -- ROS word b54
   "1000000000100000000010000011001010110011010000010111000000000101010100000000000000000100000100000000",  -- ROS word b55
   "0000000001000000000000000000000000000000000000010110101000000101101000000000000000000000000011100000",  -- ROS word b56
   "0000000001000000000000000000000000000000000000010110101000000101101000000000000000000000000011100000",  -- ROS word b57
   "0000000000100000000000000000000000001011111000010111101010000000000010000000000000000100000100000000",  -- ROS word bd4
   "0000000000000000000010000000000000000001111000010101100110000100000000000000000000000000000100000000",  -- ROS word bd5
   "0000000000100000000101010100000000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word bd6
   "0000000000100000000101010100011000000000000000000100000000000011000010000000000000000100000100000000",  -- ROS word bd7
   "1000000000010010010110000100010000000101000000011000101000000100000000000010000000000000000000110000",  -- ROS word c54
   "0000000000010010010110000100010000000101000000011000101000000100000000000010000000000000000100001000",  -- ROS word c55
   "1000000000000000000000100000000000000000000000011000100000000100000010010110100001000010000100000000",  -- ROS word c56
   "0000001010000000000000000000000000100000000000101101010010000000000000000000000000010100010100000000",  -- ROS word c57
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word cd4
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word cd5
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word cd6
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word cd7
   "1000000000000111000000000101110000000000000101011010000100000100010101001100000000000001101101001000",  -- ROS word d54
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word d55
   "1000000000000111000011000101011000000000000000011010010110000100010101001100100001000011101001001000",  -- ROS word d56
   "0000000000000111000000000101011000000000000000011010010110000100010101001100000000000011101001001000",  -- ROS word d57
   "1000000001010000000010000000000000000100100000011100100110000100000010000000000000000101011101000000",  -- ROS word dd4
   "0000000000000111100010000000000000000000000100111100100100000100000010000000000000000000110100110000",  -- ROS word dd5
   "1000000000000000000010110001001000000000000000011101000000000000000010000000000000000000110011100000",  -- ROS word dd6
   "1000001010000111000010000101101000001100100000011011001100000100000011000100000000000110000101000000",  -- ROS word dd7
   "1000000001000000000000000000000000000000000000011100100110000100000010000000000000000100000001000000",  -- ROS word e54
   "0000000000000111100010000000000000000000000100111100100100000100000010000000000000000000110100110000",  -- ROS word e55
   "1000000001000000000000110000000000000000000000011100100110000100000000000000000000000001011101000000",  -- ROS word e56
   "1001010001010000000010000000000000000100001010011101010100010100000000000000000000110001011000000000",  -- ROS word e57
   "0000001001000000000010000000000000000000000001011101101010000000000010000000000000000000000100000000",  -- ROS word ed4
   "1000000000000000010100100110101000000000000000011101100000000000000001010000100001000000000100000000",  -- ROS word ed5
   "0000000001010000010110001000000000000100011000011110001100000100000001010000100001000010000100001000",  -- ROS word ed6
   "0000000000000011100011010000000000001100111000011101100000000110001000000000000000000101101000110000",  -- ROS word ed7
   "1000000000001011100010000101101000000000000000011110101010000100000000000000000000000100000100000000",  -- ROS word f54
   "0000000000000000000010000000000000000000000100111110100010000100000000000000000000000000000100000000",  -- ROS word f55
   "1010100000000000000010000000000000000000000000011110101000000100000010000000100001000100000100000000",  -- ROS word f56
   "0100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",  -- ROS word f57
   "1011010000010111100010000000000000001011100101010110100100000000000010000000000000000100110100110000",  -- ROS word fd4
   "1000000000000111100010000110111001000000000101010110100100000100000000000000000000000100110100110000",  -- ROS word fd5
   "0000000000000111100000000110111111010000000101010110100100000100000000000000000000000100110100110000",  -- ROS word fd6
   "0000010000000000000010011000000011010000000000010111010010000100000000000000000000011000000100000000"   -- ROS word fd7
);
 
  signal addr_s : STD_LOGIC_VECTOR (0 to 11);
begin
  addr_s <= addr_i(5 to 9) & addr_i(0 to 4) & addr_i(10 to 11);
  process (clk_i)
  begin
    if (clk_i'event and clk_i = '1') then
	   if (rst='1') then
		  data_o <= (others=>'0');
		elsif (hlt='0' and hclk='1') then
  	     data_o <= ros_mem_s(to_integer(unsigned(addr_s)));
		end if;
	 end if;
  end process;
end Behavioral;

